module testModule();
    reg clk, rst;
    reg port_1;

    
    always @(posedge clk or negedge rst) begin
            
    end

    

    always @(posedge clk or negedge rst) begin
        
    end
    
endmodule //testModule
