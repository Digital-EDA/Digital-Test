#     Copyright (c) 2022 SMIC                                                       
#     Filename:      RAM64.lef                                                   
#     IP code:       S018RF2P                                                         
#     Version:       0.2.b                                                        
#     CreateDate:    Mon Oct 31 21:45:38 CST 2022                                                     
                    
#    LEF for 2-PORT Register File                                                               
#    SMIC 0.18um G Logic Process                                                       
#    Configuration: -instname RAM64 -rows 16 -bits 24 -mux 4  



# DISCLAIMER                                                                           #
#                                                                                      #  
#   SMIC hereby provides the quality information to you but makes no claims,           #
# promises or guarantees about the accuracy, completeness, or adequacy of the          #
# information herein. The information contained herein is provided on an "AS IS"       #
# basis without any warranty, and SMIC assumes no obligation to provide support        #
# of any kind or otherwise maintain the information.                                   #  
#   SMIC disclaims any representation that the information does not infringe any       #
# intellectual property rights or proprietary rights of any third parties. SMIC        #
# makes no other warranty, whether express, implied or statutory as to any             #
# matter whatsoever, including but not limited to the accuracy or sufficiency of       #
# any information or the merchantability and fitness for a particular purpose.         #
# Neither SMIC nor any of its representatives shall be liable for any cause of         #
# action incurred to connect to this service.                                          #  
#                                                                                      #
# STATEMENT OF USE AND CONFIDENTIALITY                                                 #  
#                                                                                      #  
#   The following/attached material contains confidential and proprietary              #  
# information of SMIC. This material is based upon information which SMIC              #  
# considers reliable, but SMIC neither represents nor warrants that such               #
# information is accurate or complete, and it must not be relied upon as such.         #
# This information was prepared for informational purposes and is for the use          #
# by SMIC's customer only. SMIC reserves the right to make changes in the              #  
# information at any time without notice.                                              #  
#   No part of this information may be reproduced, transmitted, transcribed,           #  
# stored in a retrieval system, or translated into any human or computer               # 
# language, in any form or by any means, electronic, mechanical, magnetic,             #  
# optical, chemical, manual, or otherwise, without the prior written consent of        #
# SMIC. Any unauthorized use or disclosure of this material is strictly                #  
# prohibited and may be unlawful. By accepting this material, the receiving            #  
# party shall be deemed to have acknowledged, accepted, and agreed to be bound         #
# by the foregoing limitations and restrictions. Thank you.                            #  
#                                                                                      #  


MACRO RAM64
CLASS BLOCK ;
ORIGIN 0 0 ;
SIZE 659.38 BY 76.2 ;
SYMMETRY X Y R90 ;

PIN QA[11]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 8.905 75.56 9.975 76.2 ;
LAYER METAL2 ;
RECT 8.905 75.56 9.975 76.2 ;
LAYER METAL3 ;
RECT 8.905 75.56 9.975 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[11]

PIN DB[11]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL2 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL3 ;
RECT 18.725 0.0 19.795 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[11]

PIN QA[10]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 32.145 75.56 33.215 76.2 ;
LAYER METAL2 ;
RECT 32.145 75.56 33.215 76.2 ;
LAYER METAL3 ;
RECT 32.145 75.56 33.215 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[10]

PIN DB[10]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL2 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL3 ;
RECT 41.965 0.0 43.035 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[10]

PIN QA[9]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 55.385 75.56 56.455 76.2 ;
LAYER METAL2 ;
RECT 55.385 75.56 56.455 76.2 ;
LAYER METAL3 ;
RECT 55.385 75.56 56.455 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[9]

PIN DB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL2 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL3 ;
RECT 65.205 0.0 66.275 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[9]

PIN QA[8]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 78.625 75.56 79.695 76.2 ;
LAYER METAL2 ;
RECT 78.625 75.56 79.695 76.2 ;
LAYER METAL3 ;
RECT 78.625 75.56 79.695 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[8]

PIN DB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL2 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL3 ;
RECT 88.445 0.0 89.515 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[8]

PIN QA[7]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 101.865 75.56 102.935 76.2 ;
LAYER METAL2 ;
RECT 101.865 75.56 102.935 76.2 ;
LAYER METAL3 ;
RECT 101.865 75.56 102.935 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[7]

PIN DB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL2 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL3 ;
RECT 111.685 0.0 112.755 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[7]

PIN QA[6]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 125.105 75.56 126.175 76.2 ;
LAYER METAL2 ;
RECT 125.105 75.56 126.175 76.2 ;
LAYER METAL3 ;
RECT 125.105 75.56 126.175 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[6]

PIN DB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL2 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL3 ;
RECT 134.925 0.0 135.995 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[6]

PIN QA[5]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 148.345 75.56 149.415 76.2 ;
LAYER METAL2 ;
RECT 148.345 75.56 149.415 76.2 ;
LAYER METAL3 ;
RECT 148.345 75.56 149.415 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[5]

PIN DB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL2 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL3 ;
RECT 158.165 0.0 159.235 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[5]

PIN QA[4]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 171.585 75.56 172.655 76.2 ;
LAYER METAL2 ;
RECT 171.585 75.56 172.655 76.2 ;
LAYER METAL3 ;
RECT 171.585 75.56 172.655 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[4]

PIN DB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL2 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL3 ;
RECT 181.405 0.0 182.475 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[4]

PIN QA[3]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 194.825 75.56 195.895 76.2 ;
LAYER METAL2 ;
RECT 194.825 75.56 195.895 76.2 ;
LAYER METAL3 ;
RECT 194.825 75.56 195.895 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[3]

PIN DB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL2 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL3 ;
RECT 204.645 0.0 205.715 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[3]

PIN QA[2]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 218.065 75.56 219.135 76.2 ;
LAYER METAL2 ;
RECT 218.065 75.56 219.135 76.2 ;
LAYER METAL3 ;
RECT 218.065 75.56 219.135 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[2]

PIN DB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL2 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL3 ;
RECT 227.885 0.0 228.955 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[2]

PIN QA[1]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 241.305 75.56 242.375 76.2 ;
LAYER METAL2 ;
RECT 241.305 75.56 242.375 76.2 ;
LAYER METAL3 ;
RECT 241.305 75.56 242.375 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[1]

PIN DB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL2 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL3 ;
RECT 251.125 0.0 252.195 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[1]

PIN QA[0]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 264.545 75.56 265.615 76.2 ;
LAYER METAL2 ;
RECT 264.545 75.56 265.615 76.2 ;
LAYER METAL3 ;
RECT 264.545 75.56 265.615 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[0]

PIN DB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL2 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL3 ;
RECT 274.365 0.0 275.435 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[0]

PIN CLKB
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL2 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL3 ;
RECT 297.105 0.0 297.605 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKB

PIN AA[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 297.655 75.56 298.905 76.2 ;
LAYER METAL2 ;
RECT 297.655 75.56 298.905 76.2 ;
LAYER METAL3 ;
RECT 297.655 75.56 298.905 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[0]

PIN AA[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 302.505 75.56 303.755 76.2 ;
LAYER METAL2 ;
RECT 302.505 75.56 303.755 76.2 ;
LAYER METAL3 ;
RECT 302.505 75.56 303.755 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[1]

PIN CENB
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL2 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL3 ;
RECT 306.72 0.0 307.22 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENB

PIN AA[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 312.875 75.56 314.525 76.2 ;
LAYER METAL2 ;
RECT 312.875 75.56 314.125 76.2 ;
LAYER METAL3 ;
RECT 312.875 75.56 314.125 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[4]

PIN AA[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 320.815 75.56 322.465 76.2 ;
LAYER METAL2 ;
RECT 320.815 75.56 322.065 76.2 ;
LAYER METAL3 ;
RECT 320.815 75.56 322.065 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[3]

PIN AB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 323.45 0.0 325.015 0.64 ;
LAYER METAL2 ;
RECT 323.765 0.0 325.015 0.64 ;
LAYER METAL3 ;
RECT 323.765 0.0 325.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[5]

PIN AA[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.755 75.56 330.405 76.2 ;
LAYER METAL2 ;
RECT 328.755 75.56 330.005 76.2 ;
LAYER METAL3 ;
RECT 328.755 75.56 330.005 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[2]

PIN AB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.975 0.0 330.625 0.64 ;
LAYER METAL2 ;
RECT 329.375 0.0 330.625 0.64 ;
LAYER METAL3 ;
RECT 329.375 0.0 330.625 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[2]

PIN AA[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.365 75.56 335.93 76.2 ;
LAYER METAL2 ;
RECT 334.365 75.56 335.615 76.2 ;
LAYER METAL3 ;
RECT 334.365 75.56 335.615 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[5]

PIN AB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 336.915 0.0 338.565 0.64 ;
LAYER METAL2 ;
RECT 337.315 0.0 338.565 0.64 ;
LAYER METAL3 ;
RECT 337.315 0.0 338.565 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[3]

PIN AB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 344.855 0.0 346.505 0.64 ;
LAYER METAL2 ;
RECT 345.255 0.0 346.505 0.64 ;
LAYER METAL3 ;
RECT 345.255 0.0 346.505 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[4]

PIN CENA
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 354.005 75.13 354.505 76.2 ;
LAYER METAL2 ;
RECT 354.005 75.13 354.505 76.2 ;
LAYER METAL3 ;
RECT 354.005 75.13 354.505 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENA

PIN AB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 355.625 0.0 356.875 0.64 ;
LAYER METAL2 ;
RECT 355.625 0.0 356.875 0.64 ;
LAYER METAL3 ;
RECT 355.625 0.0 356.875 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[1]

PIN AB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 360.475 0.0 361.725 0.64 ;
LAYER METAL2 ;
RECT 360.475 0.0 361.725 0.64 ;
LAYER METAL3 ;
RECT 360.475 0.0 361.725 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[0]

PIN CLKA
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 363.41 75.13 363.91 76.2 ;
LAYER METAL2 ;
RECT 363.41 75.13 363.91 76.2 ;
LAYER METAL3 ;
RECT 363.41 75.13 363.91 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKA

PIN DB[12]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 383.945 0.0 385.015 0.64 ;
LAYER METAL2 ;
RECT 383.945 0.0 385.015 0.64 ;
LAYER METAL3 ;
RECT 383.945 0.0 385.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[12]

PIN QA[12]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 393.765 75.56 394.835 76.2 ;
LAYER METAL2 ;
RECT 393.765 75.56 394.835 76.2 ;
LAYER METAL3 ;
RECT 393.765 75.56 394.835 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[12]

PIN DB[13]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 407.185 0.0 408.255 0.64 ;
LAYER METAL2 ;
RECT 407.185 0.0 408.255 0.64 ;
LAYER METAL3 ;
RECT 407.185 0.0 408.255 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[13]

PIN QA[13]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 417.005 75.56 418.075 76.2 ;
LAYER METAL2 ;
RECT 417.005 75.56 418.075 76.2 ;
LAYER METAL3 ;
RECT 417.005 75.56 418.075 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[13]

PIN DB[14]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 430.425 0.0 431.495 0.64 ;
LAYER METAL2 ;
RECT 430.425 0.0 431.495 0.64 ;
LAYER METAL3 ;
RECT 430.425 0.0 431.495 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[14]

PIN QA[14]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 440.245 75.56 441.315 76.2 ;
LAYER METAL2 ;
RECT 440.245 75.56 441.315 76.2 ;
LAYER METAL3 ;
RECT 440.245 75.56 441.315 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[14]

PIN DB[15]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 453.665 0.0 454.735 0.64 ;
LAYER METAL2 ;
RECT 453.665 0.0 454.735 0.64 ;
LAYER METAL3 ;
RECT 453.665 0.0 454.735 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[15]

PIN QA[15]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 463.485 75.56 464.555 76.2 ;
LAYER METAL2 ;
RECT 463.485 75.56 464.555 76.2 ;
LAYER METAL3 ;
RECT 463.485 75.56 464.555 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[15]

PIN DB[16]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 476.905 0.0 477.975 0.64 ;
LAYER METAL2 ;
RECT 476.905 0.0 477.975 0.64 ;
LAYER METAL3 ;
RECT 476.905 0.0 477.975 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[16]

PIN QA[16]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 486.725 75.56 487.795 76.2 ;
LAYER METAL2 ;
RECT 486.725 75.56 487.795 76.2 ;
LAYER METAL3 ;
RECT 486.725 75.56 487.795 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[16]

PIN DB[17]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 500.145 0.0 501.215 0.64 ;
LAYER METAL2 ;
RECT 500.145 0.0 501.215 0.64 ;
LAYER METAL3 ;
RECT 500.145 0.0 501.215 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[17]

PIN QA[17]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 509.965 75.56 511.035 76.2 ;
LAYER METAL2 ;
RECT 509.965 75.56 511.035 76.2 ;
LAYER METAL3 ;
RECT 509.965 75.56 511.035 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[17]

PIN DB[18]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 523.385 0.0 524.455 0.64 ;
LAYER METAL2 ;
RECT 523.385 0.0 524.455 0.64 ;
LAYER METAL3 ;
RECT 523.385 0.0 524.455 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[18]

PIN QA[18]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 533.205 75.56 534.275 76.2 ;
LAYER METAL2 ;
RECT 533.205 75.56 534.275 76.2 ;
LAYER METAL3 ;
RECT 533.205 75.56 534.275 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[18]

PIN DB[19]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 546.625 0.0 547.695 0.64 ;
LAYER METAL2 ;
RECT 546.625 0.0 547.695 0.64 ;
LAYER METAL3 ;
RECT 546.625 0.0 547.695 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[19]

PIN QA[19]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 556.445 75.56 557.515 76.2 ;
LAYER METAL2 ;
RECT 556.445 75.56 557.515 76.2 ;
LAYER METAL3 ;
RECT 556.445 75.56 557.515 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[19]

PIN DB[20]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 569.865 0.0 570.935 0.64 ;
LAYER METAL2 ;
RECT 569.865 0.0 570.935 0.64 ;
LAYER METAL3 ;
RECT 569.865 0.0 570.935 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[20]

PIN QA[20]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 579.685 75.56 580.755 76.2 ;
LAYER METAL2 ;
RECT 579.685 75.56 580.755 76.2 ;
LAYER METAL3 ;
RECT 579.685 75.56 580.755 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[20]

PIN DB[21]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 593.105 0.0 594.175 0.64 ;
LAYER METAL2 ;
RECT 593.105 0.0 594.175 0.64 ;
LAYER METAL3 ;
RECT 593.105 0.0 594.175 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[21]

PIN QA[21]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 602.925 75.56 603.995 76.2 ;
LAYER METAL2 ;
RECT 602.925 75.56 603.995 76.2 ;
LAYER METAL3 ;
RECT 602.925 75.56 603.995 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[21]

PIN DB[22]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 616.345 0.0 617.415 0.64 ;
LAYER METAL2 ;
RECT 616.345 0.0 617.415 0.64 ;
LAYER METAL3 ;
RECT 616.345 0.0 617.415 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[22]

PIN QA[22]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 626.165 75.56 627.235 76.2 ;
LAYER METAL2 ;
RECT 626.165 75.56 627.235 76.2 ;
LAYER METAL3 ;
RECT 626.165 75.56 627.235 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[22]

PIN DB[23]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 639.585 0.0 640.655 0.64 ;
LAYER METAL2 ;
RECT 639.585 0.0 640.655 0.64 ;
LAYER METAL3 ;
RECT 639.585 0.0 640.655 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[23]

PIN QA[23]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 649.405 75.56 650.475 76.2 ;
LAYER METAL2 ;
RECT 649.405 75.56 650.475 76.2 ;
LAYER METAL3 ;
RECT 649.405 75.56 650.475 76.2 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[23]

PIN VSS
DIRECTION INOUT ;
USE GROUND ;
PORT
LAYER METAL4 ;
RECT 279.475 0.0 283.475 76.2 ;
LAYER METAL4 ;
RECT 290.475 0.0 294.475 76.2 ;
LAYER METAL4 ;
RECT 301.475 0.0 305.475 76.2 ;
LAYER METAL4 ;
RECT 312.475 0.0 316.475 76.2 ;
LAYER METAL4 ;
RECT 323.475 0.0 327.475 76.2 ;
LAYER METAL4 ;
RECT 331.905 0.0 335.905 76.2 ;
LAYER METAL4 ;
RECT 342.905 0.0 346.905 76.2 ;
LAYER METAL4 ;
RECT 353.905 0.0 357.905 76.2 ;
LAYER METAL4 ;
RECT 364.905 0.0 368.905 76.2 ;
LAYER METAL4 ;
RECT 375.905 0.0 379.905 76.2 ;
LAYER METAL4 ;
RECT 267.855 0.0 271.855 76.2 ;
LAYER METAL4 ;
RECT 256.235 0.0 260.235 76.2 ;
LAYER METAL4 ;
RECT 244.615 0.0 248.615 76.2 ;
LAYER METAL4 ;
RECT 232.995 0.0 236.995 76.2 ;
LAYER METAL4 ;
RECT 221.375 0.0 225.375 76.2 ;
LAYER METAL4 ;
RECT 209.755 0.0 213.755 76.2 ;
LAYER METAL4 ;
RECT 198.135 0.0 202.135 76.2 ;
LAYER METAL4 ;
RECT 186.515 0.0 190.515 76.2 ;
LAYER METAL4 ;
RECT 174.895 0.0 178.895 76.2 ;
LAYER METAL4 ;
RECT 163.275 0.0 167.275 76.2 ;
LAYER METAL4 ;
RECT 151.655 0.0 155.655 76.2 ;
LAYER METAL4 ;
RECT 140.035 0.0 144.035 76.2 ;
LAYER METAL4 ;
RECT 128.415 0.0 132.415 76.2 ;
LAYER METAL4 ;
RECT 116.795 0.0 120.795 76.2 ;
LAYER METAL4 ;
RECT 105.175 0.0 109.175 76.2 ;
LAYER METAL4 ;
RECT 93.555 0.0 97.555 76.2 ;
LAYER METAL4 ;
RECT 81.935 0.0 85.935 76.2 ;
LAYER METAL4 ;
RECT 70.315 0.0 74.315 76.2 ;
LAYER METAL4 ;
RECT 58.695 0.0 62.695 76.2 ;
LAYER METAL4 ;
RECT 47.075 0.0 51.075 76.2 ;
LAYER METAL4 ;
RECT 35.455 0.0 39.455 76.2 ;
LAYER METAL4 ;
RECT 23.835 0.0 27.835 76.2 ;
LAYER METAL4 ;
RECT 12.215 0.0 16.215 76.2 ;
LAYER METAL4 ;
RECT 0.595 0.0 4.595 76.2 ;
LAYER METAL4 ;
RECT 387.525 0.0 391.525 76.2 ;
LAYER METAL4 ;
RECT 399.145 0.0 403.145 76.2 ;
LAYER METAL4 ;
RECT 410.765 0.0 414.765 76.2 ;
LAYER METAL4 ;
RECT 422.385 0.0 426.385 76.2 ;
LAYER METAL4 ;
RECT 434.005 0.0 438.005 76.2 ;
LAYER METAL4 ;
RECT 445.625 0.0 449.625 76.2 ;
LAYER METAL4 ;
RECT 457.245 0.0 461.245 76.2 ;
LAYER METAL4 ;
RECT 468.865 0.0 472.865 76.2 ;
LAYER METAL4 ;
RECT 480.485 0.0 484.485 76.2 ;
LAYER METAL4 ;
RECT 492.105 0.0 496.105 76.2 ;
LAYER METAL4 ;
RECT 503.725 0.0 507.725 76.2 ;
LAYER METAL4 ;
RECT 515.345 0.0 519.345 76.2 ;
LAYER METAL4 ;
RECT 526.965 0.0 530.965 76.2 ;
LAYER METAL4 ;
RECT 538.585 0.0 542.585 76.2 ;
LAYER METAL4 ;
RECT 550.205 0.0 554.205 76.2 ;
LAYER METAL4 ;
RECT 561.825 0.0 565.825 76.2 ;
LAYER METAL4 ;
RECT 573.445 0.0 577.445 76.2 ;
LAYER METAL4 ;
RECT 585.065 0.0 589.065 76.2 ;
LAYER METAL4 ;
RECT 596.685 0.0 600.685 76.2 ;
LAYER METAL4 ;
RECT 608.305 0.0 612.305 76.2 ;
LAYER METAL4 ;
RECT 619.925 0.0 623.925 76.2 ;
LAYER METAL4 ;
RECT 631.545 0.0 635.545 76.2 ;
LAYER METAL4 ;
RECT 643.165 0.0 647.165 76.2 ;
LAYER METAL4 ;
RECT 654.785 0.0 658.785 76.2 ;
END
END VSS

PIN VDD
DIRECTION INOUT ;
USE POWER ;
PORT
LAYER METAL4 ;
RECT 284.975 0.0 288.975 76.2 ;
LAYER METAL4 ;
RECT 295.975 0.0 299.975 76.2 ;
LAYER METAL4 ;
RECT 306.975 0.0 310.975 76.2 ;
LAYER METAL4 ;
RECT 317.975 0.0 321.975 76.2 ;
LAYER METAL4 ;
RECT 337.405 0.0 341.405 76.2 ;
LAYER METAL4 ;
RECT 348.405 0.0 352.405 76.2 ;
LAYER METAL4 ;
RECT 359.405 0.0 363.405 76.2 ;
LAYER METAL4 ;
RECT 370.405 0.0 374.405 76.2 ;
LAYER METAL4 ;
RECT 273.665 0.0 277.665 76.2 ;
LAYER METAL4 ;
RECT 262.045 0.0 266.045 76.2 ;
LAYER METAL4 ;
RECT 250.425 0.0 254.425 76.2 ;
LAYER METAL4 ;
RECT 238.805 0.0 242.805 76.2 ;
LAYER METAL4 ;
RECT 227.185 0.0 231.185 76.2 ;
LAYER METAL4 ;
RECT 215.565 0.0 219.565 76.2 ;
LAYER METAL4 ;
RECT 203.945 0.0 207.945 76.2 ;
LAYER METAL4 ;
RECT 192.325 0.0 196.325 76.2 ;
LAYER METAL4 ;
RECT 180.705 0.0 184.705 76.2 ;
LAYER METAL4 ;
RECT 169.085 0.0 173.085 76.2 ;
LAYER METAL4 ;
RECT 157.465 0.0 161.465 76.2 ;
LAYER METAL4 ;
RECT 145.845 0.0 149.845 76.2 ;
LAYER METAL4 ;
RECT 134.225 0.0 138.225 76.2 ;
LAYER METAL4 ;
RECT 122.605 0.0 126.605 76.2 ;
LAYER METAL4 ;
RECT 110.985 0.0 114.985 76.2 ;
LAYER METAL4 ;
RECT 99.365 0.0 103.365 76.2 ;
LAYER METAL4 ;
RECT 87.745 0.0 91.745 76.2 ;
LAYER METAL4 ;
RECT 76.125 0.0 80.125 76.2 ;
LAYER METAL4 ;
RECT 64.505 0.0 68.505 76.2 ;
LAYER METAL4 ;
RECT 52.885 0.0 56.885 76.2 ;
LAYER METAL4 ;
RECT 41.265 0.0 45.265 76.2 ;
LAYER METAL4 ;
RECT 29.645 0.0 33.645 76.2 ;
LAYER METAL4 ;
RECT 18.025 0.0 22.025 76.2 ;
LAYER METAL4 ;
RECT 6.405 0.0 10.405 76.2 ;
LAYER METAL4 ;
RECT 381.715 0.0 385.715 76.2 ;
LAYER METAL4 ;
RECT 393.335 0.0 397.335 76.2 ;
LAYER METAL4 ;
RECT 404.955 0.0 408.955 76.2 ;
LAYER METAL4 ;
RECT 416.575 0.0 420.575 76.2 ;
LAYER METAL4 ;
RECT 428.195 0.0 432.195 76.2 ;
LAYER METAL4 ;
RECT 439.815 0.0 443.815 76.2 ;
LAYER METAL4 ;
RECT 451.435 0.0 455.435 76.2 ;
LAYER METAL4 ;
RECT 463.055 0.0 467.055 76.2 ;
LAYER METAL4 ;
RECT 474.675 0.0 478.675 76.2 ;
LAYER METAL4 ;
RECT 486.295 0.0 490.295 76.2 ;
LAYER METAL4 ;
RECT 497.915 0.0 501.915 76.2 ;
LAYER METAL4 ;
RECT 509.535 0.0 513.535 76.2 ;
LAYER METAL4 ;
RECT 521.155 0.0 525.155 76.2 ;
LAYER METAL4 ;
RECT 532.775 0.0 536.775 76.2 ;
LAYER METAL4 ;
RECT 544.395 0.0 548.395 76.2 ;
LAYER METAL4 ;
RECT 556.015 0.0 560.015 76.2 ;
LAYER METAL4 ;
RECT 567.635 0.0 571.635 76.2 ;
LAYER METAL4 ;
RECT 579.255 0.0 583.255 76.2 ;
LAYER METAL4 ;
RECT 590.875 0.0 594.875 76.2 ;
LAYER METAL4 ;
RECT 602.495 0.0 606.495 76.2 ;
LAYER METAL4 ;
RECT 614.115 0.0 618.115 76.2 ;
LAYER METAL4 ;
RECT 625.735 0.0 629.735 76.2 ;
LAYER METAL4 ;
RECT 637.355 0.0 641.355 76.2 ;
LAYER METAL4 ;
RECT 648.975 0.0 652.975 76.2 ;
END
END VDD

OBS
LAYER VIA12 ;
RECT  0.000 0.000 659.380 76.200 ;
LAYER VIA23 ;
RECT  0.000 0.000 659.380 76.200 ;
LAYER VIA34 ;
RECT  0.000 0.000 659.380 76.200 ;
LAYER METAL1 ;
POLYGON 0.000 0.000 18.495 0.000 18.495 0.870 20.025 0.870 20.025 0.000
 41.735 0.000 41.735 0.870 43.265 0.870 43.265 0.000 64.975 0.000
 64.975 0.870 66.505 0.870 66.505 0.000 88.215 0.000 88.215 0.870
 89.745 0.870 89.745 0.000 111.455 0.000 111.455 0.870 112.985 0.870
 112.985 0.000 134.695 0.000 134.695 0.870 136.225 0.870 136.225 0.000
 157.935 0.000 157.935 0.870 159.465 0.870 159.465 0.000 181.175 0.000
 181.175 0.870 182.705 0.870 182.705 0.000 204.415 0.000 204.415 0.870
 205.945 0.870 205.945 0.000 227.655 0.000 227.655 0.870 229.185 0.870
 229.185 0.000 250.895 0.000 250.895 0.870 252.425 0.870 252.425 0.000
 274.135 0.000 274.135 0.870 275.665 0.870 275.665 0.000 296.875 0.000
 296.875 1.300 297.835 1.300 297.835 0.000 306.490 0.000 306.490 1.300
 307.450 1.300 307.450 0.000 323.220 0.000 323.220 0.870 325.245 0.870
 325.245 0.000 328.745 0.000 328.745 0.870 330.855 0.870 330.855 0.000
 336.685 0.000 336.685 0.870 338.795 0.870 338.795 0.000 344.625 0.000
 344.625 0.870 346.735 0.870 346.735 0.000 355.395 0.000 355.395 0.870
 357.105 0.870 357.105 0.000 360.245 0.000 360.245 0.870 361.955 0.870
 361.955 0.000 383.715 0.000 383.715 0.870 385.245 0.870 385.245 0.000
 406.955 0.000 406.955 0.870 408.485 0.870 408.485 0.000 430.195 0.000
 430.195 0.870 431.725 0.870 431.725 0.000 453.435 0.000 453.435 0.870
 454.965 0.870 454.965 0.000 476.675 0.000 476.675 0.870 478.205 0.870
 478.205 0.000 499.915 0.000 499.915 0.870 501.445 0.870 501.445 0.000
 523.155 0.000 523.155 0.870 524.685 0.870 524.685 0.000 546.395 0.000
 546.395 0.870 547.925 0.870 547.925 0.000 569.635 0.000 569.635 0.870
 571.165 0.870 571.165 0.000 592.875 0.000 592.875 0.870 594.405 0.870
 594.405 0.000 616.115 0.000 616.115 0.870 617.645 0.870 617.645 0.000
 639.355 0.000 639.355 0.870 640.885 0.870 640.885 0.000 659.380 0.000
 659.380 76.200 650.705 76.200 650.705 75.330 649.175 75.330 649.175 76.200
 627.465 76.200 627.465 75.330 625.935 75.330 625.935 76.200 604.225 76.200
 604.225 75.330 602.695 75.330 602.695 76.200 580.985 76.200 580.985 75.330
 579.455 75.330 579.455 76.200 557.745 76.200 557.745 75.330 556.215 75.330
 556.215 76.200 534.505 76.200 534.505 75.330 532.975 75.330 532.975 76.200
 511.265 76.200 511.265 75.330 509.735 75.330 509.735 76.200 488.025 76.200
 488.025 75.330 486.495 75.330 486.495 76.200 464.785 76.200 464.785 75.330
 463.255 75.330 463.255 76.200 441.545 76.200 441.545 75.330 440.015 75.330
 440.015 76.200 418.305 76.200 418.305 75.330 416.775 75.330 416.775 76.200
 395.065 76.200 395.065 75.330 393.535 75.330 393.535 76.200 364.140 76.200
 364.140 74.900 363.180 74.900 363.180 76.200 354.735 76.200 354.735 74.900
 353.775 74.900 353.775 76.200 336.160 76.200 336.160 75.330 334.135 75.330
 334.135 76.200 330.635 76.200 330.635 75.330 328.525 75.330 328.525 76.200
 322.695 76.200 322.695 75.330 320.585 75.330 320.585 76.200 314.755 76.200
 314.755 75.330 312.645 75.330 312.645 76.200 303.985 76.200 303.985 75.330
 302.275 75.330 302.275 76.200 299.135 76.200 299.135 75.330 297.425 75.330
 297.425 76.200 265.845 76.200 265.845 75.330 264.315 75.330 264.315 76.200
 242.605 76.200 242.605 75.330 241.075 75.330 241.075 76.200 219.365 76.200
 219.365 75.330 217.835 75.330 217.835 76.200 196.125 76.200 196.125 75.330
 194.595 75.330 194.595 76.200 172.885 76.200 172.885 75.330 171.355 75.330
 171.355 76.200 149.645 76.200 149.645 75.330 148.115 75.330 148.115 76.200
 126.405 76.200 126.405 75.330 124.875 75.330 124.875 76.200 103.165 76.200
 103.165 75.330 101.635 75.330 101.635 76.200 79.925 76.200 79.925 75.330
 78.395 75.330 78.395 76.200 56.685 76.200 56.685 75.330 55.155 75.330
 55.155 76.200 33.445 76.200 33.445 75.330 31.915 75.330 31.915 76.200
 10.205 76.200 10.205 75.330 8.675 75.330 8.675 76.200 0.000 76.200
 ;
LAYER METAL2 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.095 0.000 329.095 0.920 330.905 0.920 330.905 0.000
 337.035 0.000 337.035 0.920 338.845 0.920 338.845 0.000 344.975 0.000
 344.975 0.920 346.785 0.920 346.785 0.000 355.345 0.000 355.345 0.920
 357.155 0.920 357.155 0.000 360.195 0.000 360.195 0.920 362.005 0.920
 362.005 0.000 383.665 0.000 383.665 0.920 385.295 0.920 385.295 0.000
 406.905 0.000 406.905 0.920 408.535 0.920 408.535 0.000 430.145 0.000
 430.145 0.920 431.775 0.920 431.775 0.000 453.385 0.000 453.385 0.920
 455.015 0.920 455.015 0.000 476.625 0.000 476.625 0.920 478.255 0.920
 478.255 0.000 499.865 0.000 499.865 0.920 501.495 0.920 501.495 0.000
 523.105 0.000 523.105 0.920 524.735 0.920 524.735 0.000 546.345 0.000
 546.345 0.920 547.975 0.920 547.975 0.000 569.585 0.000 569.585 0.920
 571.215 0.920 571.215 0.000 592.825 0.000 592.825 0.920 594.455 0.920
 594.455 0.000 616.065 0.000 616.065 0.920 617.695 0.920 617.695 0.000
 639.305 0.000 639.305 0.920 640.935 0.920 640.935 0.000 659.380 0.000
 659.380 76.200 650.755 76.200 650.755 75.280 649.125 75.280 649.125 76.200
 627.515 76.200 627.515 75.280 625.885 75.280 625.885 76.200 604.275 76.200
 604.275 75.280 602.645 75.280 602.645 76.200 581.035 76.200 581.035 75.280
 579.405 75.280 579.405 76.200 557.795 76.200 557.795 75.280 556.165 75.280
 556.165 76.200 534.555 76.200 534.555 75.280 532.925 75.280 532.925 76.200
 511.315 76.200 511.315 75.280 509.685 75.280 509.685 76.200 488.075 76.200
 488.075 75.280 486.445 75.280 486.445 76.200 464.835 76.200 464.835 75.280
 463.205 75.280 463.205 76.200 441.595 76.200 441.595 75.280 439.965 75.280
 439.965 76.200 418.355 76.200 418.355 75.280 416.725 75.280 416.725 76.200
 395.115 76.200 395.115 75.280 393.485 75.280 393.485 76.200 364.190 76.200
 364.190 74.850 363.130 74.850 363.130 76.200 354.785 76.200 354.785 74.850
 353.725 74.850 353.725 76.200 335.895 76.200 335.895 75.280 334.085 75.280
 334.085 76.200 330.285 76.200 330.285 75.280 328.475 75.280 328.475 76.200
 322.345 76.200 322.345 75.280 320.535 75.280 320.535 76.200 314.405 76.200
 314.405 75.280 312.595 75.280 312.595 76.200 304.035 76.200 304.035 75.280
 302.225 75.280 302.225 76.200 299.185 76.200 299.185 75.280 297.375 75.280
 297.375 76.200 265.895 76.200 265.895 75.280 264.265 75.280 264.265 76.200
 242.655 76.200 242.655 75.280 241.025 75.280 241.025 76.200 219.415 76.200
 219.415 75.280 217.785 75.280 217.785 76.200 196.175 76.200 196.175 75.280
 194.545 75.280 194.545 76.200 172.935 76.200 172.935 75.280 171.305 75.280
 171.305 76.200 149.695 76.200 149.695 75.280 148.065 75.280 148.065 76.200
 126.455 76.200 126.455 75.280 124.825 75.280 124.825 76.200 103.215 76.200
 103.215 75.280 101.585 75.280 101.585 76.200 79.975 76.200 79.975 75.280
 78.345 75.280 78.345 76.200 56.735 76.200 56.735 75.280 55.105 75.280
 55.105 76.200 33.495 76.200 33.495 75.280 31.865 75.280 31.865 76.200
 10.255 76.200 10.255 75.280 8.625 75.280 8.625 76.200 0.000 76.200
 ;
LAYER METAL3 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.095 0.000 329.095 0.920 330.905 0.920 330.905 0.000
 337.035 0.000 337.035 0.920 338.845 0.920 338.845 0.000 344.975 0.000
 344.975 0.920 346.785 0.920 346.785 0.000 355.345 0.000 355.345 0.920
 357.155 0.920 357.155 0.000 360.195 0.000 360.195 0.920 362.005 0.920
 362.005 0.000 383.665 0.000 383.665 0.920 385.295 0.920 385.295 0.000
 406.905 0.000 406.905 0.920 408.535 0.920 408.535 0.000 430.145 0.000
 430.145 0.920 431.775 0.920 431.775 0.000 453.385 0.000 453.385 0.920
 455.015 0.920 455.015 0.000 476.625 0.000 476.625 0.920 478.255 0.920
 478.255 0.000 499.865 0.000 499.865 0.920 501.495 0.920 501.495 0.000
 523.105 0.000 523.105 0.920 524.735 0.920 524.735 0.000 546.345 0.000
 546.345 0.920 547.975 0.920 547.975 0.000 569.585 0.000 569.585 0.920
 571.215 0.920 571.215 0.000 592.825 0.000 592.825 0.920 594.455 0.920
 594.455 0.000 616.065 0.000 616.065 0.920 617.695 0.920 617.695 0.000
 639.305 0.000 639.305 0.920 640.935 0.920 640.935 0.000 659.380 0.000
 659.380 76.200 650.755 76.200 650.755 75.280 649.125 75.280 649.125 76.200
 627.515 76.200 627.515 75.280 625.885 75.280 625.885 76.200 604.275 76.200
 604.275 75.280 602.645 75.280 602.645 76.200 581.035 76.200 581.035 75.280
 579.405 75.280 579.405 76.200 557.795 76.200 557.795 75.280 556.165 75.280
 556.165 76.200 534.555 76.200 534.555 75.280 532.925 75.280 532.925 76.200
 511.315 76.200 511.315 75.280 509.685 75.280 509.685 76.200 488.075 76.200
 488.075 75.280 486.445 75.280 486.445 76.200 464.835 76.200 464.835 75.280
 463.205 75.280 463.205 76.200 441.595 76.200 441.595 75.280 439.965 75.280
 439.965 76.200 418.355 76.200 418.355 75.280 416.725 75.280 416.725 76.200
 395.115 76.200 395.115 75.280 393.485 75.280 393.485 76.200 364.190 76.200
 364.190 74.850 363.130 74.850 363.130 76.200 354.785 76.200 354.785 74.850
 353.725 74.850 353.725 76.200 335.895 76.200 335.895 75.280 334.085 75.280
 334.085 76.200 330.285 76.200 330.285 75.280 328.475 75.280 328.475 76.200
 322.345 76.200 322.345 75.280 320.535 75.280 320.535 76.200 314.405 76.200
 314.405 75.280 312.595 75.280 312.595 76.200 304.035 76.200 304.035 75.280
 302.225 75.280 302.225 76.200 299.185 76.200 299.185 75.280 297.375 75.280
 297.375 76.200 265.895 76.200 265.895 75.280 264.265 75.280 264.265 76.200
 242.655 76.200 242.655 75.280 241.025 75.280 241.025 76.200 219.415 76.200
 219.415 75.280 217.785 75.280 217.785 76.200 196.175 76.200 196.175 75.280
 194.545 75.280 194.545 76.200 172.935 76.200 172.935 75.280 171.305 75.280
 171.305 76.200 149.695 76.200 149.695 75.280 148.065 75.280 148.065 76.200
 126.455 76.200 126.455 75.280 124.825 75.280 124.825 76.200 103.215 76.200
 103.215 75.280 101.585 75.280 101.585 76.200 79.975 76.200 79.975 75.280
 78.345 75.280 78.345 76.200 56.735 76.200 56.735 75.280 55.105 75.280
 55.105 76.200 33.495 76.200 33.495 75.280 31.865 75.280 31.865 76.200
 10.255 76.200 10.255 75.280 8.625 75.280 8.625 76.200 0.000 76.200
 ;
END
END RAM64
END LIBRARY
