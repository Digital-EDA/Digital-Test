#     Copyright (c) 2022 SMIC                                                       
#     Filename:      RAM256.lef                                                   
#     IP code:       S018RF2P                                                         
#     Version:       0.2.b                                                        
#     CreateDate:    Mon Oct 31 21:43:58 CST 2022                                                     
                    
#    LEF for 2-PORT Register File                                                               
#    SMIC 0.18um G Logic Process                                                       
#    Configuration: -instname RAM256 -rows 64 -bits 24 -mux 4  



# DISCLAIMER                                                                           #
#                                                                                      #  
#   SMIC hereby provides the quality information to you but makes no claims,           #
# promises or guarantees about the accuracy, completeness, or adequacy of the          #
# information herein. The information contained herein is provided on an "AS IS"       #
# basis without any warranty, and SMIC assumes no obligation to provide support        #
# of any kind or otherwise maintain the information.                                   #  
#   SMIC disclaims any representation that the information does not infringe any       #
# intellectual property rights or proprietary rights of any third parties. SMIC        #
# makes no other warranty, whether express, implied or statutory as to any             #
# matter whatsoever, including but not limited to the accuracy or sufficiency of       #
# any information or the merchantability and fitness for a particular purpose.         #
# Neither SMIC nor any of its representatives shall be liable for any cause of         #
# action incurred to connect to this service.                                          #  
#                                                                                      #
# STATEMENT OF USE AND CONFIDENTIALITY                                                 #  
#                                                                                      #  
#   The following/attached material contains confidential and proprietary              #  
# information of SMIC. This material is based upon information which SMIC              #  
# considers reliable, but SMIC neither represents nor warrants that such               #
# information is accurate or complete, and it must not be relied upon as such.         #
# This information was prepared for informational purposes and is for the use          #
# by SMIC's customer only. SMIC reserves the right to make changes in the              #  
# information at any time without notice.                                              #  
#   No part of this information may be reproduced, transmitted, transcribed,           #  
# stored in a retrieval system, or translated into any human or computer               # 
# language, in any form or by any means, electronic, mechanical, magnetic,             #  
# optical, chemical, manual, or otherwise, without the prior written consent of        #
# SMIC. Any unauthorized use or disclosure of this material is strictly                #  
# prohibited and may be unlawful. By accepting this material, the receiving            #  
# party shall be deemed to have acknowledged, accepted, and agreed to be bound         #
# by the foregoing limitations and restrictions. Thank you.                            #  
#                                                                                      #  


MACRO RAM256
CLASS BLOCK ;
ORIGIN 0 0 ;
SIZE 670.9 BY 159.945 ;
SYMMETRY X Y R90 ;

PIN QA[11]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 8.905 159.305 9.975 159.945 ;
LAYER METAL2 ;
RECT 8.905 159.305 9.975 159.945 ;
LAYER METAL3 ;
RECT 8.905 159.305 9.975 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[11]

PIN DB[11]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL2 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL3 ;
RECT 18.725 0.0 19.795 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[11]

PIN QA[10]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 32.145 159.305 33.215 159.945 ;
LAYER METAL2 ;
RECT 32.145 159.305 33.215 159.945 ;
LAYER METAL3 ;
RECT 32.145 159.305 33.215 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[10]

PIN DB[10]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL2 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL3 ;
RECT 41.965 0.0 43.035 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[10]

PIN QA[9]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 55.385 159.305 56.455 159.945 ;
LAYER METAL2 ;
RECT 55.385 159.305 56.455 159.945 ;
LAYER METAL3 ;
RECT 55.385 159.305 56.455 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[9]

PIN DB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL2 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL3 ;
RECT 65.205 0.0 66.275 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[9]

PIN QA[8]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 78.625 159.305 79.695 159.945 ;
LAYER METAL2 ;
RECT 78.625 159.305 79.695 159.945 ;
LAYER METAL3 ;
RECT 78.625 159.305 79.695 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[8]

PIN DB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL2 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL3 ;
RECT 88.445 0.0 89.515 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[8]

PIN QA[7]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 101.865 159.305 102.935 159.945 ;
LAYER METAL2 ;
RECT 101.865 159.305 102.935 159.945 ;
LAYER METAL3 ;
RECT 101.865 159.305 102.935 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[7]

PIN DB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL2 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL3 ;
RECT 111.685 0.0 112.755 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[7]

PIN QA[6]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 125.105 159.305 126.175 159.945 ;
LAYER METAL2 ;
RECT 125.105 159.305 126.175 159.945 ;
LAYER METAL3 ;
RECT 125.105 159.305 126.175 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[6]

PIN DB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL2 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL3 ;
RECT 134.925 0.0 135.995 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[6]

PIN QA[5]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 148.345 159.305 149.415 159.945 ;
LAYER METAL2 ;
RECT 148.345 159.305 149.415 159.945 ;
LAYER METAL3 ;
RECT 148.345 159.305 149.415 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[5]

PIN DB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL2 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL3 ;
RECT 158.165 0.0 159.235 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[5]

PIN QA[4]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 171.585 159.305 172.655 159.945 ;
LAYER METAL2 ;
RECT 171.585 159.305 172.655 159.945 ;
LAYER METAL3 ;
RECT 171.585 159.305 172.655 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[4]

PIN DB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL2 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL3 ;
RECT 181.405 0.0 182.475 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[4]

PIN QA[3]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 194.825 159.305 195.895 159.945 ;
LAYER METAL2 ;
RECT 194.825 159.305 195.895 159.945 ;
LAYER METAL3 ;
RECT 194.825 159.305 195.895 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[3]

PIN DB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL2 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL3 ;
RECT 204.645 0.0 205.715 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[3]

PIN QA[2]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 218.065 159.305 219.135 159.945 ;
LAYER METAL2 ;
RECT 218.065 159.305 219.135 159.945 ;
LAYER METAL3 ;
RECT 218.065 159.305 219.135 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[2]

PIN DB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL2 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL3 ;
RECT 227.885 0.0 228.955 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[2]

PIN QA[1]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 241.305 159.305 242.375 159.945 ;
LAYER METAL2 ;
RECT 241.305 159.305 242.375 159.945 ;
LAYER METAL3 ;
RECT 241.305 159.305 242.375 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[1]

PIN DB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL2 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL3 ;
RECT 251.125 0.0 252.195 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[1]

PIN QA[0]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 264.545 159.305 265.615 159.945 ;
LAYER METAL2 ;
RECT 264.545 159.305 265.615 159.945 ;
LAYER METAL3 ;
RECT 264.545 159.305 265.615 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[0]

PIN DB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL2 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL3 ;
RECT 274.365 0.0 275.435 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[0]

PIN CLKB
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL2 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL3 ;
RECT 297.105 0.0 297.605 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKB

PIN AA[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 297.655 159.305 298.905 159.945 ;
LAYER METAL2 ;
RECT 297.655 159.305 298.905 159.945 ;
LAYER METAL3 ;
RECT 297.655 159.305 298.905 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[0]

PIN AA[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 302.505 159.305 303.755 159.945 ;
LAYER METAL2 ;
RECT 302.505 159.305 303.755 159.945 ;
LAYER METAL3 ;
RECT 302.505 159.305 303.755 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[1]

PIN CENB
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL2 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL3 ;
RECT 306.72 0.0 307.22 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENB

PIN AA[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 312.875 159.305 314.525 159.945 ;
LAYER METAL2 ;
RECT 312.875 159.305 314.125 159.945 ;
LAYER METAL3 ;
RECT 312.875 159.305 314.125 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[4]

PIN AA[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 320.815 159.305 322.465 159.945 ;
LAYER METAL2 ;
RECT 320.815 159.305 322.065 159.945 ;
LAYER METAL3 ;
RECT 320.815 159.305 322.065 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[3]

PIN AB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 323.45 0.0 325.015 0.64 ;
LAYER METAL2 ;
RECT 323.765 0.0 325.015 0.64 ;
LAYER METAL3 ;
RECT 323.765 0.0 325.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[7]

PIN AA[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.755 159.305 330.405 159.945 ;
LAYER METAL2 ;
RECT 328.755 159.305 330.005 159.945 ;
LAYER METAL3 ;
RECT 328.755 159.305 330.005 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[2]

PIN AB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 329.21 0.0 330.775 0.64 ;
LAYER METAL2 ;
RECT 329.525 0.0 330.775 0.64 ;
LAYER METAL3 ;
RECT 329.525 0.0 330.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[6]

PIN AA[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.365 159.305 335.93 159.945 ;
LAYER METAL2 ;
RECT 334.365 159.305 335.615 159.945 ;
LAYER METAL3 ;
RECT 334.365 159.305 335.615 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[5]

PIN AB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.97 0.0 336.535 0.64 ;
LAYER METAL2 ;
RECT 335.285 0.0 336.535 0.64 ;
LAYER METAL3 ;
RECT 335.285 0.0 336.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[5]

PIN AA[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.125 159.305 341.69 159.945 ;
LAYER METAL2 ;
RECT 340.125 159.305 341.375 159.945 ;
LAYER METAL3 ;
RECT 340.125 159.305 341.375 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[6]

PIN AB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.495 0.0 342.145 0.64 ;
LAYER METAL2 ;
RECT 340.895 0.0 342.145 0.64 ;
LAYER METAL3 ;
RECT 340.895 0.0 342.145 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[2]

PIN AA[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 345.885 159.305 347.45 159.945 ;
LAYER METAL2 ;
RECT 345.885 159.305 347.135 159.945 ;
LAYER METAL3 ;
RECT 345.885 159.305 347.135 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[7]

PIN AB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 348.435 0.0 350.085 0.64 ;
LAYER METAL2 ;
RECT 348.835 0.0 350.085 0.64 ;
LAYER METAL3 ;
RECT 348.835 0.0 350.085 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[3]

PIN AB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 356.375 0.0 358.025 0.64 ;
LAYER METAL2 ;
RECT 356.775 0.0 358.025 0.64 ;
LAYER METAL3 ;
RECT 356.775 0.0 358.025 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[4]

PIN CENA
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 365.525 158.875 366.025 159.945 ;
LAYER METAL2 ;
RECT 365.525 158.875 366.025 159.945 ;
LAYER METAL3 ;
RECT 365.525 158.875 366.025 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENA

PIN AB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 367.145 0.0 368.395 0.64 ;
LAYER METAL2 ;
RECT 367.145 0.0 368.395 0.64 ;
LAYER METAL3 ;
RECT 367.145 0.0 368.395 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[1]

PIN AB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 371.995 0.0 373.245 0.64 ;
LAYER METAL2 ;
RECT 371.995 0.0 373.245 0.64 ;
LAYER METAL3 ;
RECT 371.995 0.0 373.245 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[0]

PIN CLKA
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 374.93 158.875 375.43 159.945 ;
LAYER METAL2 ;
RECT 374.93 158.875 375.43 159.945 ;
LAYER METAL3 ;
RECT 374.93 158.875 375.43 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKA

PIN DB[12]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 395.465 0.0 396.535 0.64 ;
LAYER METAL2 ;
RECT 395.465 0.0 396.535 0.64 ;
LAYER METAL3 ;
RECT 395.465 0.0 396.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[12]

PIN QA[12]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 405.285 159.305 406.355 159.945 ;
LAYER METAL2 ;
RECT 405.285 159.305 406.355 159.945 ;
LAYER METAL3 ;
RECT 405.285 159.305 406.355 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[12]

PIN DB[13]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 418.705 0.0 419.775 0.64 ;
LAYER METAL2 ;
RECT 418.705 0.0 419.775 0.64 ;
LAYER METAL3 ;
RECT 418.705 0.0 419.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[13]

PIN QA[13]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 428.525 159.305 429.595 159.945 ;
LAYER METAL2 ;
RECT 428.525 159.305 429.595 159.945 ;
LAYER METAL3 ;
RECT 428.525 159.305 429.595 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[13]

PIN DB[14]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 441.945 0.0 443.015 0.64 ;
LAYER METAL2 ;
RECT 441.945 0.0 443.015 0.64 ;
LAYER METAL3 ;
RECT 441.945 0.0 443.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[14]

PIN QA[14]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 451.765 159.305 452.835 159.945 ;
LAYER METAL2 ;
RECT 451.765 159.305 452.835 159.945 ;
LAYER METAL3 ;
RECT 451.765 159.305 452.835 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[14]

PIN DB[15]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 465.185 0.0 466.255 0.64 ;
LAYER METAL2 ;
RECT 465.185 0.0 466.255 0.64 ;
LAYER METAL3 ;
RECT 465.185 0.0 466.255 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[15]

PIN QA[15]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 475.005 159.305 476.075 159.945 ;
LAYER METAL2 ;
RECT 475.005 159.305 476.075 159.945 ;
LAYER METAL3 ;
RECT 475.005 159.305 476.075 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[15]

PIN DB[16]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 488.425 0.0 489.495 0.64 ;
LAYER METAL2 ;
RECT 488.425 0.0 489.495 0.64 ;
LAYER METAL3 ;
RECT 488.425 0.0 489.495 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[16]

PIN QA[16]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 498.245 159.305 499.315 159.945 ;
LAYER METAL2 ;
RECT 498.245 159.305 499.315 159.945 ;
LAYER METAL3 ;
RECT 498.245 159.305 499.315 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[16]

PIN DB[17]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 511.665 0.0 512.735 0.64 ;
LAYER METAL2 ;
RECT 511.665 0.0 512.735 0.64 ;
LAYER METAL3 ;
RECT 511.665 0.0 512.735 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[17]

PIN QA[17]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 521.485 159.305 522.555 159.945 ;
LAYER METAL2 ;
RECT 521.485 159.305 522.555 159.945 ;
LAYER METAL3 ;
RECT 521.485 159.305 522.555 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[17]

PIN DB[18]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 534.905 0.0 535.975 0.64 ;
LAYER METAL2 ;
RECT 534.905 0.0 535.975 0.64 ;
LAYER METAL3 ;
RECT 534.905 0.0 535.975 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[18]

PIN QA[18]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 544.725 159.305 545.795 159.945 ;
LAYER METAL2 ;
RECT 544.725 159.305 545.795 159.945 ;
LAYER METAL3 ;
RECT 544.725 159.305 545.795 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[18]

PIN DB[19]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 558.145 0.0 559.215 0.64 ;
LAYER METAL2 ;
RECT 558.145 0.0 559.215 0.64 ;
LAYER METAL3 ;
RECT 558.145 0.0 559.215 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[19]

PIN QA[19]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 567.965 159.305 569.035 159.945 ;
LAYER METAL2 ;
RECT 567.965 159.305 569.035 159.945 ;
LAYER METAL3 ;
RECT 567.965 159.305 569.035 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[19]

PIN DB[20]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 581.385 0.0 582.455 0.64 ;
LAYER METAL2 ;
RECT 581.385 0.0 582.455 0.64 ;
LAYER METAL3 ;
RECT 581.385 0.0 582.455 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[20]

PIN QA[20]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 591.205 159.305 592.275 159.945 ;
LAYER METAL2 ;
RECT 591.205 159.305 592.275 159.945 ;
LAYER METAL3 ;
RECT 591.205 159.305 592.275 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[20]

PIN DB[21]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 604.625 0.0 605.695 0.64 ;
LAYER METAL2 ;
RECT 604.625 0.0 605.695 0.64 ;
LAYER METAL3 ;
RECT 604.625 0.0 605.695 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[21]

PIN QA[21]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 614.445 159.305 615.515 159.945 ;
LAYER METAL2 ;
RECT 614.445 159.305 615.515 159.945 ;
LAYER METAL3 ;
RECT 614.445 159.305 615.515 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[21]

PIN DB[22]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 627.865 0.0 628.935 0.64 ;
LAYER METAL2 ;
RECT 627.865 0.0 628.935 0.64 ;
LAYER METAL3 ;
RECT 627.865 0.0 628.935 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[22]

PIN QA[22]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 637.685 159.305 638.755 159.945 ;
LAYER METAL2 ;
RECT 637.685 159.305 638.755 159.945 ;
LAYER METAL3 ;
RECT 637.685 159.305 638.755 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[22]

PIN DB[23]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 651.105 0.0 652.175 0.64 ;
LAYER METAL2 ;
RECT 651.105 0.0 652.175 0.64 ;
LAYER METAL3 ;
RECT 651.105 0.0 652.175 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[23]

PIN QA[23]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 660.925 159.305 661.995 159.945 ;
LAYER METAL2 ;
RECT 660.925 159.305 661.995 159.945 ;
LAYER METAL3 ;
RECT 660.925 159.305 661.995 159.945 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[23]

PIN VSS
DIRECTION INOUT ;
USE GROUND ;
PORT
LAYER METAL4 ;
RECT 279.475 0.0 283.475 159.945 ;
LAYER METAL4 ;
RECT 290.475 0.0 294.475 159.945 ;
LAYER METAL4 ;
RECT 301.475 0.0 305.475 159.945 ;
LAYER METAL4 ;
RECT 312.475 0.0 316.475 159.945 ;
LAYER METAL4 ;
RECT 323.475 0.0 327.475 159.945 ;
LAYER METAL4 ;
RECT 343.425 0.0 347.425 159.945 ;
LAYER METAL4 ;
RECT 354.425 0.0 358.425 159.945 ;
LAYER METAL4 ;
RECT 365.425 0.0 369.425 159.945 ;
LAYER METAL4 ;
RECT 376.425 0.0 380.425 159.945 ;
LAYER METAL4 ;
RECT 387.425 0.0 391.425 159.945 ;
LAYER METAL4 ;
RECT 267.855 0.0 271.855 159.945 ;
LAYER METAL4 ;
RECT 256.235 0.0 260.235 159.945 ;
LAYER METAL4 ;
RECT 244.615 0.0 248.615 159.945 ;
LAYER METAL4 ;
RECT 232.995 0.0 236.995 159.945 ;
LAYER METAL4 ;
RECT 221.375 0.0 225.375 159.945 ;
LAYER METAL4 ;
RECT 209.755 0.0 213.755 159.945 ;
LAYER METAL4 ;
RECT 198.135 0.0 202.135 159.945 ;
LAYER METAL4 ;
RECT 186.515 0.0 190.515 159.945 ;
LAYER METAL4 ;
RECT 174.895 0.0 178.895 159.945 ;
LAYER METAL4 ;
RECT 163.275 0.0 167.275 159.945 ;
LAYER METAL4 ;
RECT 151.655 0.0 155.655 159.945 ;
LAYER METAL4 ;
RECT 140.035 0.0 144.035 159.945 ;
LAYER METAL4 ;
RECT 128.415 0.0 132.415 159.945 ;
LAYER METAL4 ;
RECT 116.795 0.0 120.795 159.945 ;
LAYER METAL4 ;
RECT 105.175 0.0 109.175 159.945 ;
LAYER METAL4 ;
RECT 93.555 0.0 97.555 159.945 ;
LAYER METAL4 ;
RECT 81.935 0.0 85.935 159.945 ;
LAYER METAL4 ;
RECT 70.315 0.0 74.315 159.945 ;
LAYER METAL4 ;
RECT 58.695 0.0 62.695 159.945 ;
LAYER METAL4 ;
RECT 47.075 0.0 51.075 159.945 ;
LAYER METAL4 ;
RECT 35.455 0.0 39.455 159.945 ;
LAYER METAL4 ;
RECT 23.835 0.0 27.835 159.945 ;
LAYER METAL4 ;
RECT 12.215 0.0 16.215 159.945 ;
LAYER METAL4 ;
RECT 0.595 0.0 4.595 159.945 ;
LAYER METAL4 ;
RECT 399.045 0.0 403.045 159.945 ;
LAYER METAL4 ;
RECT 410.665 0.0 414.665 159.945 ;
LAYER METAL4 ;
RECT 422.285 0.0 426.285 159.945 ;
LAYER METAL4 ;
RECT 433.905 0.0 437.905 159.945 ;
LAYER METAL4 ;
RECT 445.525 0.0 449.525 159.945 ;
LAYER METAL4 ;
RECT 457.145 0.0 461.145 159.945 ;
LAYER METAL4 ;
RECT 468.765 0.0 472.765 159.945 ;
LAYER METAL4 ;
RECT 480.385 0.0 484.385 159.945 ;
LAYER METAL4 ;
RECT 492.005 0.0 496.005 159.945 ;
LAYER METAL4 ;
RECT 503.625 0.0 507.625 159.945 ;
LAYER METAL4 ;
RECT 515.245 0.0 519.245 159.945 ;
LAYER METAL4 ;
RECT 526.865 0.0 530.865 159.945 ;
LAYER METAL4 ;
RECT 538.485 0.0 542.485 159.945 ;
LAYER METAL4 ;
RECT 550.105 0.0 554.105 159.945 ;
LAYER METAL4 ;
RECT 561.725 0.0 565.725 159.945 ;
LAYER METAL4 ;
RECT 573.345 0.0 577.345 159.945 ;
LAYER METAL4 ;
RECT 584.965 0.0 588.965 159.945 ;
LAYER METAL4 ;
RECT 596.585 0.0 600.585 159.945 ;
LAYER METAL4 ;
RECT 608.205 0.0 612.205 159.945 ;
LAYER METAL4 ;
RECT 619.825 0.0 623.825 159.945 ;
LAYER METAL4 ;
RECT 631.445 0.0 635.445 159.945 ;
LAYER METAL4 ;
RECT 643.065 0.0 647.065 159.945 ;
LAYER METAL4 ;
RECT 654.685 0.0 658.685 159.945 ;
LAYER METAL4 ;
RECT 666.305 0.0 670.305 159.945 ;
END
END VSS

PIN VDD
DIRECTION INOUT ;
USE POWER ;
PORT
LAYER METAL4 ;
RECT 284.975 0.0 288.975 159.945 ;
LAYER METAL4 ;
RECT 295.975 0.0 299.975 159.945 ;
LAYER METAL4 ;
RECT 306.975 0.0 310.975 159.945 ;
LAYER METAL4 ;
RECT 317.975 0.0 321.975 159.945 ;
LAYER METAL4 ;
RECT 328.975 0.0 332.975 159.945 ;
LAYER METAL4 ;
RECT 337.925 0.0 341.925 159.945 ;
LAYER METAL4 ;
RECT 348.925 0.0 352.925 159.945 ;
LAYER METAL4 ;
RECT 359.925 0.0 363.925 159.945 ;
LAYER METAL4 ;
RECT 370.925 0.0 374.925 159.945 ;
LAYER METAL4 ;
RECT 381.925 0.0 385.925 159.945 ;
LAYER METAL4 ;
RECT 273.665 0.0 277.665 159.945 ;
LAYER METAL4 ;
RECT 262.045 0.0 266.045 159.945 ;
LAYER METAL4 ;
RECT 250.425 0.0 254.425 159.945 ;
LAYER METAL4 ;
RECT 238.805 0.0 242.805 159.945 ;
LAYER METAL4 ;
RECT 227.185 0.0 231.185 159.945 ;
LAYER METAL4 ;
RECT 215.565 0.0 219.565 159.945 ;
LAYER METAL4 ;
RECT 203.945 0.0 207.945 159.945 ;
LAYER METAL4 ;
RECT 192.325 0.0 196.325 159.945 ;
LAYER METAL4 ;
RECT 180.705 0.0 184.705 159.945 ;
LAYER METAL4 ;
RECT 169.085 0.0 173.085 159.945 ;
LAYER METAL4 ;
RECT 157.465 0.0 161.465 159.945 ;
LAYER METAL4 ;
RECT 145.845 0.0 149.845 159.945 ;
LAYER METAL4 ;
RECT 134.225 0.0 138.225 159.945 ;
LAYER METAL4 ;
RECT 122.605 0.0 126.605 159.945 ;
LAYER METAL4 ;
RECT 110.985 0.0 114.985 159.945 ;
LAYER METAL4 ;
RECT 99.365 0.0 103.365 159.945 ;
LAYER METAL4 ;
RECT 87.745 0.0 91.745 159.945 ;
LAYER METAL4 ;
RECT 76.125 0.0 80.125 159.945 ;
LAYER METAL4 ;
RECT 64.505 0.0 68.505 159.945 ;
LAYER METAL4 ;
RECT 52.885 0.0 56.885 159.945 ;
LAYER METAL4 ;
RECT 41.265 0.0 45.265 159.945 ;
LAYER METAL4 ;
RECT 29.645 0.0 33.645 159.945 ;
LAYER METAL4 ;
RECT 18.025 0.0 22.025 159.945 ;
LAYER METAL4 ;
RECT 6.405 0.0 10.405 159.945 ;
LAYER METAL4 ;
RECT 393.235 0.0 397.235 159.945 ;
LAYER METAL4 ;
RECT 404.855 0.0 408.855 159.945 ;
LAYER METAL4 ;
RECT 416.475 0.0 420.475 159.945 ;
LAYER METAL4 ;
RECT 428.095 0.0 432.095 159.945 ;
LAYER METAL4 ;
RECT 439.715 0.0 443.715 159.945 ;
LAYER METAL4 ;
RECT 451.335 0.0 455.335 159.945 ;
LAYER METAL4 ;
RECT 462.955 0.0 466.955 159.945 ;
LAYER METAL4 ;
RECT 474.575 0.0 478.575 159.945 ;
LAYER METAL4 ;
RECT 486.195 0.0 490.195 159.945 ;
LAYER METAL4 ;
RECT 497.815 0.0 501.815 159.945 ;
LAYER METAL4 ;
RECT 509.435 0.0 513.435 159.945 ;
LAYER METAL4 ;
RECT 521.055 0.0 525.055 159.945 ;
LAYER METAL4 ;
RECT 532.675 0.0 536.675 159.945 ;
LAYER METAL4 ;
RECT 544.295 0.0 548.295 159.945 ;
LAYER METAL4 ;
RECT 555.915 0.0 559.915 159.945 ;
LAYER METAL4 ;
RECT 567.535 0.0 571.535 159.945 ;
LAYER METAL4 ;
RECT 579.155 0.0 583.155 159.945 ;
LAYER METAL4 ;
RECT 590.775 0.0 594.775 159.945 ;
LAYER METAL4 ;
RECT 602.395 0.0 606.395 159.945 ;
LAYER METAL4 ;
RECT 614.015 0.0 618.015 159.945 ;
LAYER METAL4 ;
RECT 625.635 0.0 629.635 159.945 ;
LAYER METAL4 ;
RECT 637.255 0.0 641.255 159.945 ;
LAYER METAL4 ;
RECT 648.875 0.0 652.875 159.945 ;
LAYER METAL4 ;
RECT 660.495 0.0 664.495 159.945 ;
END
END VDD

OBS
LAYER VIA12 ;
RECT  0.000 0.000 670.900 159.945 ;
LAYER VIA23 ;
RECT  0.000 0.000 670.900 159.945 ;
LAYER VIA34 ;
RECT  0.000 0.000 670.900 159.945 ;
LAYER METAL1 ;
POLYGON 0.000 0.000 18.495 0.000 18.495 0.870 20.025 0.870 20.025 0.000
 41.735 0.000 41.735 0.870 43.265 0.870 43.265 0.000 64.975 0.000
 64.975 0.870 66.505 0.870 66.505 0.000 88.215 0.000 88.215 0.870
 89.745 0.870 89.745 0.000 111.455 0.000 111.455 0.870 112.985 0.870
 112.985 0.000 134.695 0.000 134.695 0.870 136.225 0.870 136.225 0.000
 157.935 0.000 157.935 0.870 159.465 0.870 159.465 0.000 181.175 0.000
 181.175 0.870 182.705 0.870 182.705 0.000 204.415 0.000 204.415 0.870
 205.945 0.870 205.945 0.000 227.655 0.000 227.655 0.870 229.185 0.870
 229.185 0.000 250.895 0.000 250.895 0.870 252.425 0.870 252.425 0.000
 274.135 0.000 274.135 0.870 275.665 0.870 275.665 0.000 296.875 0.000
 296.875 1.300 297.835 1.300 297.835 0.000 306.490 0.000 306.490 1.300
 307.450 1.300 307.450 0.000 323.220 0.000 323.220 0.870 325.245 0.870
 325.245 0.000 328.980 0.000 328.980 0.870 331.005 0.870 331.005 0.000
 334.740 0.000 334.740 0.870 336.765 0.870 336.765 0.000 340.265 0.000
 340.265 0.870 342.375 0.870 342.375 0.000 348.205 0.000 348.205 0.870
 350.315 0.870 350.315 0.000 356.145 0.000 356.145 0.870 358.255 0.870
 358.255 0.000 366.915 0.000 366.915 0.870 368.625 0.870 368.625 0.000
 371.765 0.000 371.765 0.870 373.475 0.870 373.475 0.000 395.235 0.000
 395.235 0.870 396.765 0.870 396.765 0.000 418.475 0.000 418.475 0.870
 420.005 0.870 420.005 0.000 441.715 0.000 441.715 0.870 443.245 0.870
 443.245 0.000 464.955 0.000 464.955 0.870 466.485 0.870 466.485 0.000
 488.195 0.000 488.195 0.870 489.725 0.870 489.725 0.000 511.435 0.000
 511.435 0.870 512.965 0.870 512.965 0.000 534.675 0.000 534.675 0.870
 536.205 0.870 536.205 0.000 557.915 0.000 557.915 0.870 559.445 0.870
 559.445 0.000 581.155 0.000 581.155 0.870 582.685 0.870 582.685 0.000
 604.395 0.000 604.395 0.870 605.925 0.870 605.925 0.000 627.635 0.000
 627.635 0.870 629.165 0.870 629.165 0.000 650.875 0.000 650.875 0.870
 652.405 0.870 652.405 0.000 670.900 0.000 670.900 159.945 662.225 159.945 662.225 159.075 660.695 159.075 660.695 159.945
 638.985 159.945 638.985 159.075 637.455 159.075 637.455 159.945 615.745 159.945
 615.745 159.075 614.215 159.075 614.215 159.945 592.505 159.945 592.505 159.075
 590.975 159.075 590.975 159.945 569.265 159.945 569.265 159.075 567.735 159.075
 567.735 159.945 546.025 159.945 546.025 159.075 544.495 159.075 544.495 159.945
 522.785 159.945 522.785 159.075 521.255 159.075 521.255 159.945 499.545 159.945
 499.545 159.075 498.015 159.075 498.015 159.945 476.305 159.945 476.305 159.075
 474.775 159.075 474.775 159.945 453.065 159.945 453.065 159.075 451.535 159.075
 451.535 159.945 429.825 159.945 429.825 159.075 428.295 159.075 428.295 159.945
 406.585 159.945 406.585 159.075 405.055 159.075 405.055 159.945 375.660 159.945
 375.660 158.645 374.700 158.645 374.700 159.945 366.255 159.945 366.255 158.645
 365.295 158.645 365.295 159.945 347.680 159.945 347.680 159.075 345.655 159.075
 345.655 159.945 341.920 159.945 341.920 159.075 339.895 159.075 339.895 159.945
 336.160 159.945 336.160 159.075 334.135 159.075 334.135 159.945 330.635 159.945
 330.635 159.075 328.525 159.075 328.525 159.945 322.695 159.945 322.695 159.075
 320.585 159.075 320.585 159.945 314.755 159.945 314.755 159.075 312.645 159.075
 312.645 159.945 303.985 159.945 303.985 159.075 302.275 159.075 302.275 159.945
 299.135 159.945 299.135 159.075 297.425 159.075 297.425 159.945 265.845 159.945
 265.845 159.075 264.315 159.075 264.315 159.945 242.605 159.945 242.605 159.075
 241.075 159.075 241.075 159.945 219.365 159.945 219.365 159.075 217.835 159.075
 217.835 159.945 196.125 159.945 196.125 159.075 194.595 159.075 194.595 159.945
 172.885 159.945 172.885 159.075 171.355 159.075 171.355 159.945 149.645 159.945
 149.645 159.075 148.115 159.075 148.115 159.945 126.405 159.945 126.405 159.075
 124.875 159.075 124.875 159.945 103.165 159.945 103.165 159.075 101.635 159.075
 101.635 159.945 79.925 159.945 79.925 159.075 78.395 159.075 78.395 159.945
 56.685 159.945 56.685 159.075 55.155 159.075 55.155 159.945 33.445 159.945
 33.445 159.075 31.915 159.075 31.915 159.945 10.205 159.945 10.205 159.075
 8.675 159.075 8.675 159.945 0.000 159.945 ;
LAYER METAL2 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 335.005 0.000 335.005 0.920 336.815 0.920 336.815 0.000 340.615 0.000
 340.615 0.920 342.425 0.920 342.425 0.000 348.555 0.000 348.555 0.920
 350.365 0.920 350.365 0.000 356.495 0.000 356.495 0.920 358.305 0.920
 358.305 0.000 366.865 0.000 366.865 0.920 368.675 0.920 368.675 0.000
 371.715 0.000 371.715 0.920 373.525 0.920 373.525 0.000 395.185 0.000
 395.185 0.920 396.815 0.920 396.815 0.000 418.425 0.000 418.425 0.920
 420.055 0.920 420.055 0.000 441.665 0.000 441.665 0.920 443.295 0.920
 443.295 0.000 464.905 0.000 464.905 0.920 466.535 0.920 466.535 0.000
 488.145 0.000 488.145 0.920 489.775 0.920 489.775 0.000 511.385 0.000
 511.385 0.920 513.015 0.920 513.015 0.000 534.625 0.000 534.625 0.920
 536.255 0.920 536.255 0.000 557.865 0.000 557.865 0.920 559.495 0.920
 559.495 0.000 581.105 0.000 581.105 0.920 582.735 0.920 582.735 0.000
 604.345 0.000 604.345 0.920 605.975 0.920 605.975 0.000 627.585 0.000
 627.585 0.920 629.215 0.920 629.215 0.000 650.825 0.000 650.825 0.920
 652.455 0.920 652.455 0.000 670.900 0.000 670.900 159.945 662.275 159.945 662.275 159.025 660.645 159.025 660.645 159.945
 639.035 159.945 639.035 159.025 637.405 159.025 637.405 159.945 615.795 159.945
 615.795 159.025 614.165 159.025 614.165 159.945 592.555 159.945 592.555 159.025
 590.925 159.025 590.925 159.945 569.315 159.945 569.315 159.025 567.685 159.025
 567.685 159.945 546.075 159.945 546.075 159.025 544.445 159.025 544.445 159.945
 522.835 159.945 522.835 159.025 521.205 159.025 521.205 159.945 499.595 159.945
 499.595 159.025 497.965 159.025 497.965 159.945 476.355 159.945 476.355 159.025
 474.725 159.025 474.725 159.945 453.115 159.945 453.115 159.025 451.485 159.025
 451.485 159.945 429.875 159.945 429.875 159.025 428.245 159.025 428.245 159.945
 406.635 159.945 406.635 159.025 405.005 159.025 405.005 159.945 375.710 159.945
 375.710 158.595 374.650 158.595 374.650 159.945 366.305 159.945 366.305 158.595
 365.245 158.595 365.245 159.945 347.415 159.945 347.415 159.025 345.605 159.025
 345.605 159.945 341.655 159.945 341.655 159.025 339.845 159.025 339.845 159.945
 335.895 159.945 335.895 159.025 334.085 159.025 334.085 159.945 330.285 159.945
 330.285 159.025 328.475 159.025 328.475 159.945 322.345 159.945 322.345 159.025
 320.535 159.025 320.535 159.945 314.405 159.945 314.405 159.025 312.595 159.025
 312.595 159.945 304.035 159.945 304.035 159.025 302.225 159.025 302.225 159.945
 299.185 159.945 299.185 159.025 297.375 159.025 297.375 159.945 265.895 159.945
 265.895 159.025 264.265 159.025 264.265 159.945 242.655 159.945 242.655 159.025
 241.025 159.025 241.025 159.945 219.415 159.945 219.415 159.025 217.785 159.025
 217.785 159.945 196.175 159.945 196.175 159.025 194.545 159.025 194.545 159.945
 172.935 159.945 172.935 159.025 171.305 159.025 171.305 159.945 149.695 159.945
 149.695 159.025 148.065 159.025 148.065 159.945 126.455 159.945 126.455 159.025
 124.825 159.025 124.825 159.945 103.215 159.945 103.215 159.025 101.585 159.025
 101.585 159.945 79.975 159.945 79.975 159.025 78.345 159.025 78.345 159.945
 56.735 159.945 56.735 159.025 55.105 159.025 55.105 159.945 33.495 159.945
 33.495 159.025 31.865 159.025 31.865 159.945 10.255 159.945 10.255 159.025
 8.625 159.025 8.625 159.945 0.000 159.945 ;
LAYER METAL3 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 335.005 0.000 335.005 0.920 336.815 0.920 336.815 0.000 340.615 0.000
 340.615 0.920 342.425 0.920 342.425 0.000 348.555 0.000 348.555 0.920
 350.365 0.920 350.365 0.000 356.495 0.000 356.495 0.920 358.305 0.920
 358.305 0.000 366.865 0.000 366.865 0.920 368.675 0.920 368.675 0.000
 371.715 0.000 371.715 0.920 373.525 0.920 373.525 0.000 395.185 0.000
 395.185 0.920 396.815 0.920 396.815 0.000 418.425 0.000 418.425 0.920
 420.055 0.920 420.055 0.000 441.665 0.000 441.665 0.920 443.295 0.920
 443.295 0.000 464.905 0.000 464.905 0.920 466.535 0.920 466.535 0.000
 488.145 0.000 488.145 0.920 489.775 0.920 489.775 0.000 511.385 0.000
 511.385 0.920 513.015 0.920 513.015 0.000 534.625 0.000 534.625 0.920
 536.255 0.920 536.255 0.000 557.865 0.000 557.865 0.920 559.495 0.920
 559.495 0.000 581.105 0.000 581.105 0.920 582.735 0.920 582.735 0.000
 604.345 0.000 604.345 0.920 605.975 0.920 605.975 0.000 627.585 0.000
 627.585 0.920 629.215 0.920 629.215 0.000 650.825 0.000 650.825 0.920
 652.455 0.920 652.455 0.000 670.900 0.000 670.900 159.945 662.275 159.945 662.275 159.025 660.645 159.025 660.645 159.945
 639.035 159.945 639.035 159.025 637.405 159.025 637.405 159.945 615.795 159.945
 615.795 159.025 614.165 159.025 614.165 159.945 592.555 159.945 592.555 159.025
 590.925 159.025 590.925 159.945 569.315 159.945 569.315 159.025 567.685 159.025
 567.685 159.945 546.075 159.945 546.075 159.025 544.445 159.025 544.445 159.945
 522.835 159.945 522.835 159.025 521.205 159.025 521.205 159.945 499.595 159.945
 499.595 159.025 497.965 159.025 497.965 159.945 476.355 159.945 476.355 159.025
 474.725 159.025 474.725 159.945 453.115 159.945 453.115 159.025 451.485 159.025
 451.485 159.945 429.875 159.945 429.875 159.025 428.245 159.025 428.245 159.945
 406.635 159.945 406.635 159.025 405.005 159.025 405.005 159.945 375.710 159.945
 375.710 158.595 374.650 158.595 374.650 159.945 366.305 159.945 366.305 158.595
 365.245 158.595 365.245 159.945 347.415 159.945 347.415 159.025 345.605 159.025
 345.605 159.945 341.655 159.945 341.655 159.025 339.845 159.025 339.845 159.945
 335.895 159.945 335.895 159.025 334.085 159.025 334.085 159.945 330.285 159.945
 330.285 159.025 328.475 159.025 328.475 159.945 322.345 159.945 322.345 159.025
 320.535 159.025 320.535 159.945 314.405 159.945 314.405 159.025 312.595 159.025
 312.595 159.945 304.035 159.945 304.035 159.025 302.225 159.025 302.225 159.945
 299.185 159.945 299.185 159.025 297.375 159.025 297.375 159.945 265.895 159.945
 265.895 159.025 264.265 159.025 264.265 159.945 242.655 159.945 242.655 159.025
 241.025 159.025 241.025 159.945 219.415 159.945 219.415 159.025 217.785 159.025
 217.785 159.945 196.175 159.945 196.175 159.025 194.545 159.025 194.545 159.945
 172.935 159.945 172.935 159.025 171.305 159.025 171.305 159.945 149.695 159.945
 149.695 159.025 148.065 159.025 148.065 159.945 126.455 159.945 126.455 159.025
 124.825 159.025 124.825 159.945 103.215 159.945 103.215 159.025 101.585 159.025
 101.585 159.945 79.975 159.945 79.975 159.025 78.345 159.025 78.345 159.945
 56.735 159.945 56.735 159.025 55.105 159.025 55.105 159.945 33.495 159.945
 33.495 159.025 31.865 159.025 31.865 159.945 10.255 159.945 10.255 159.025
 8.625 159.025 8.625 159.945 0.000 159.945 ;
END
END RAM256
END LIBRARY
