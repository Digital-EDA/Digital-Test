#     Copyright (c) 2022 SMIC                                                       
#     Filename:      RAM1024.lef                                                   
#     IP code:       S018RF2P                                                         
#     Version:       0.2.b                                                        
#     CreateDate:    Sun Sep 11 16:38:48 CST 2022                                                     
                    
#    LEF for 2-PORT Register File                                                               
#    SMIC 0.18um G Logic Process                                                       
#    Configuration: -instname RAM1024 -rows 256 -bits 24 -mux 4  



# DISCLAIMER                                                                           #
#                                                                                      #  
#   SMIC hereby provides the quality information to you but makes no claims,           #
# promises or guarantees about the accuracy, completeness, or adequacy of the          #
# information herein. The information contained herein is provided on an "AS IS"       #
# basis without any warranty, and SMIC assumes no obligation to provide support        #
# of any kind or otherwise maintain the information.                                   #  
#   SMIC disclaims any representation that the information does not infringe any       #
# intellectual property rights or proprietary rights of any third parties. SMIC        #
# makes no other warranty, whether express, implied or statutory as to any             #
# matter whatsoever, including but not limited to the accuracy or sufficiency of       #
# any information or the merchantability and fitness for a particular purpose.         #
# Neither SMIC nor any of its representatives shall be liable for any cause of         #
# action incurred to connect to this service.                                          #  
#                                                                                      #
# STATEMENT OF USE AND CONFIDENTIALITY                                                 #  
#                                                                                      #  
#   The following/attached material contains confidential and proprietary              #  
# information of SMIC. This material is based upon information which SMIC              #  
# considers reliable, but SMIC neither represents nor warrants that such               #
# information is accurate or complete, and it must not be relied upon as such.         #
# This information was prepared for informational purposes and is for the use          #
# by SMIC's customer only. SMIC reserves the right to make changes in the              #  
# information at any time without notice.                                              #  
#   No part of this information may be reproduced, transmitted, transcribed,           #  
# stored in a retrieval system, or translated into any human or computer               # 
# language, in any form or by any means, electronic, mechanical, magnetic,             #  
# optical, chemical, manual, or otherwise, without the prior written consent of        #
# SMIC. Any unauthorized use or disclosure of this material is strictly                #  
# prohibited and may be unlawful. By accepting this material, the receiving            #  
# party shall be deemed to have acknowledged, accepted, and agreed to be bound         #
# by the foregoing limitations and restrictions. Thank you.                            #  
#                                                                                      #  


MACRO RAM1024
CLASS BLOCK ;
ORIGIN 0 0 ;
SIZE 682.42 BY 496.905 ;
SYMMETRY X Y R90 ;

PIN QA[11]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 8.905 496.265 9.975 496.905 ;
LAYER METAL2 ;
RECT 8.905 496.265 9.975 496.905 ;
LAYER METAL3 ;
RECT 8.905 496.265 9.975 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[11]

PIN DB[11]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL2 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL3 ;
RECT 18.725 0.0 19.795 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[11]

PIN QA[10]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 32.145 496.265 33.215 496.905 ;
LAYER METAL2 ;
RECT 32.145 496.265 33.215 496.905 ;
LAYER METAL3 ;
RECT 32.145 496.265 33.215 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[10]

PIN DB[10]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL2 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL3 ;
RECT 41.965 0.0 43.035 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[10]

PIN QA[9]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 55.385 496.265 56.455 496.905 ;
LAYER METAL2 ;
RECT 55.385 496.265 56.455 496.905 ;
LAYER METAL3 ;
RECT 55.385 496.265 56.455 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[9]

PIN DB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL2 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL3 ;
RECT 65.205 0.0 66.275 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[9]

PIN QA[8]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 78.625 496.265 79.695 496.905 ;
LAYER METAL2 ;
RECT 78.625 496.265 79.695 496.905 ;
LAYER METAL3 ;
RECT 78.625 496.265 79.695 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[8]

PIN DB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL2 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL3 ;
RECT 88.445 0.0 89.515 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[8]

PIN QA[7]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 101.865 496.265 102.935 496.905 ;
LAYER METAL2 ;
RECT 101.865 496.265 102.935 496.905 ;
LAYER METAL3 ;
RECT 101.865 496.265 102.935 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[7]

PIN DB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL2 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL3 ;
RECT 111.685 0.0 112.755 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[7]

PIN QA[6]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 125.105 496.265 126.175 496.905 ;
LAYER METAL2 ;
RECT 125.105 496.265 126.175 496.905 ;
LAYER METAL3 ;
RECT 125.105 496.265 126.175 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[6]

PIN DB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL2 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL3 ;
RECT 134.925 0.0 135.995 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[6]

PIN QA[5]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 148.345 496.265 149.415 496.905 ;
LAYER METAL2 ;
RECT 148.345 496.265 149.415 496.905 ;
LAYER METAL3 ;
RECT 148.345 496.265 149.415 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[5]

PIN DB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL2 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL3 ;
RECT 158.165 0.0 159.235 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[5]

PIN QA[4]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 171.585 496.265 172.655 496.905 ;
LAYER METAL2 ;
RECT 171.585 496.265 172.655 496.905 ;
LAYER METAL3 ;
RECT 171.585 496.265 172.655 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[4]

PIN DB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL2 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL3 ;
RECT 181.405 0.0 182.475 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[4]

PIN QA[3]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 194.825 496.265 195.895 496.905 ;
LAYER METAL2 ;
RECT 194.825 496.265 195.895 496.905 ;
LAYER METAL3 ;
RECT 194.825 496.265 195.895 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[3]

PIN DB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL2 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL3 ;
RECT 204.645 0.0 205.715 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[3]

PIN QA[2]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 218.065 496.265 219.135 496.905 ;
LAYER METAL2 ;
RECT 218.065 496.265 219.135 496.905 ;
LAYER METAL3 ;
RECT 218.065 496.265 219.135 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[2]

PIN DB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL2 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL3 ;
RECT 227.885 0.0 228.955 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[2]

PIN QA[1]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 241.305 496.265 242.375 496.905 ;
LAYER METAL2 ;
RECT 241.305 496.265 242.375 496.905 ;
LAYER METAL3 ;
RECT 241.305 496.265 242.375 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[1]

PIN DB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL2 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL3 ;
RECT 251.125 0.0 252.195 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[1]

PIN QA[0]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 264.545 496.265 265.615 496.905 ;
LAYER METAL2 ;
RECT 264.545 496.265 265.615 496.905 ;
LAYER METAL3 ;
RECT 264.545 496.265 265.615 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[0]

PIN DB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL2 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL3 ;
RECT 274.365 0.0 275.435 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[0]

PIN CLKB
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL2 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL3 ;
RECT 297.105 0.0 297.605 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKB

PIN AA[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 297.655 496.265 298.905 496.905 ;
LAYER METAL2 ;
RECT 297.655 496.265 298.905 496.905 ;
LAYER METAL3 ;
RECT 297.655 496.265 298.905 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[0]

PIN AA[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 302.505 496.265 303.755 496.905 ;
LAYER METAL2 ;
RECT 302.505 496.265 303.755 496.905 ;
LAYER METAL3 ;
RECT 302.505 496.265 303.755 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[1]

PIN CENB
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL2 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL3 ;
RECT 306.72 0.0 307.22 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENB

PIN AA[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 312.875 496.265 314.525 496.905 ;
LAYER METAL2 ;
RECT 312.875 496.265 314.125 496.905 ;
LAYER METAL3 ;
RECT 312.875 496.265 314.125 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[4]

PIN AA[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 320.815 496.265 322.465 496.905 ;
LAYER METAL2 ;
RECT 320.815 496.265 322.065 496.905 ;
LAYER METAL3 ;
RECT 320.815 496.265 322.065 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[3]

PIN AB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 323.45 0.0 325.015 0.64 ;
LAYER METAL2 ;
RECT 323.765 0.0 325.015 0.64 ;
LAYER METAL3 ;
RECT 323.765 0.0 325.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[9]

PIN AA[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.755 496.265 330.405 496.905 ;
LAYER METAL2 ;
RECT 328.755 496.265 330.005 496.905 ;
LAYER METAL3 ;
RECT 328.755 496.265 330.005 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[2]

PIN AB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 329.21 0.0 330.775 0.64 ;
LAYER METAL2 ;
RECT 329.525 0.0 330.775 0.64 ;
LAYER METAL3 ;
RECT 329.525 0.0 330.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[8]

PIN AA[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.365 496.265 335.93 496.905 ;
LAYER METAL2 ;
RECT 334.365 496.265 335.615 496.905 ;
LAYER METAL3 ;
RECT 334.365 496.265 335.615 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[5]

PIN AB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.97 0.0 336.535 0.64 ;
LAYER METAL2 ;
RECT 335.285 0.0 336.535 0.64 ;
LAYER METAL3 ;
RECT 335.285 0.0 336.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[7]

PIN AA[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.125 496.265 341.69 496.905 ;
LAYER METAL2 ;
RECT 340.125 496.265 341.375 496.905 ;
LAYER METAL3 ;
RECT 340.125 496.265 341.375 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[6]

PIN AB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.73 0.0 342.295 0.64 ;
LAYER METAL2 ;
RECT 341.045 0.0 342.295 0.64 ;
LAYER METAL3 ;
RECT 341.045 0.0 342.295 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[6]

PIN AA[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 345.885 496.265 347.45 496.905 ;
LAYER METAL2 ;
RECT 345.885 496.265 347.135 496.905 ;
LAYER METAL3 ;
RECT 345.885 496.265 347.135 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[7]

PIN AB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 346.49 0.0 348.055 0.64 ;
LAYER METAL2 ;
RECT 346.805 0.0 348.055 0.64 ;
LAYER METAL3 ;
RECT 346.805 0.0 348.055 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[5]

PIN AA[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 351.645 496.265 353.21 496.905 ;
LAYER METAL2 ;
RECT 351.645 496.265 352.895 496.905 ;
LAYER METAL3 ;
RECT 351.645 496.265 352.895 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[8]

PIN AB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 352.015 0.0 353.665 0.64 ;
LAYER METAL2 ;
RECT 352.415 0.0 353.665 0.64 ;
LAYER METAL3 ;
RECT 352.415 0.0 353.665 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[2]

PIN AA[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 357.405 496.265 358.97 496.905 ;
LAYER METAL2 ;
RECT 357.405 496.265 358.655 496.905 ;
LAYER METAL3 ;
RECT 357.405 496.265 358.655 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[9]

PIN AB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 359.955 0.0 361.605 0.64 ;
LAYER METAL2 ;
RECT 360.355 0.0 361.605 0.64 ;
LAYER METAL3 ;
RECT 360.355 0.0 361.605 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[3]

PIN AB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 367.895 0.0 369.545 0.64 ;
LAYER METAL2 ;
RECT 368.295 0.0 369.545 0.64 ;
LAYER METAL3 ;
RECT 368.295 0.0 369.545 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[4]

PIN CENA
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 377.045 495.835 377.545 496.905 ;
LAYER METAL2 ;
RECT 377.045 495.835 377.545 496.905 ;
LAYER METAL3 ;
RECT 377.045 495.835 377.545 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENA

PIN AB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 378.665 0.0 379.915 0.64 ;
LAYER METAL2 ;
RECT 378.665 0.0 379.915 0.64 ;
LAYER METAL3 ;
RECT 378.665 0.0 379.915 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[1]

PIN AB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 383.515 0.0 384.765 0.64 ;
LAYER METAL2 ;
RECT 383.515 0.0 384.765 0.64 ;
LAYER METAL3 ;
RECT 383.515 0.0 384.765 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[0]

PIN CLKA
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 386.45 495.835 386.95 496.905 ;
LAYER METAL2 ;
RECT 386.45 495.835 386.95 496.905 ;
LAYER METAL3 ;
RECT 386.45 495.835 386.95 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKA

PIN DB[12]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 406.985 0.0 408.055 0.64 ;
LAYER METAL2 ;
RECT 406.985 0.0 408.055 0.64 ;
LAYER METAL3 ;
RECT 406.985 0.0 408.055 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[12]

PIN QA[12]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 416.805 496.265 417.875 496.905 ;
LAYER METAL2 ;
RECT 416.805 496.265 417.875 496.905 ;
LAYER METAL3 ;
RECT 416.805 496.265 417.875 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[12]

PIN DB[13]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 430.225 0.0 431.295 0.64 ;
LAYER METAL2 ;
RECT 430.225 0.0 431.295 0.64 ;
LAYER METAL3 ;
RECT 430.225 0.0 431.295 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[13]

PIN QA[13]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 440.045 496.265 441.115 496.905 ;
LAYER METAL2 ;
RECT 440.045 496.265 441.115 496.905 ;
LAYER METAL3 ;
RECT 440.045 496.265 441.115 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[13]

PIN DB[14]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 453.465 0.0 454.535 0.64 ;
LAYER METAL2 ;
RECT 453.465 0.0 454.535 0.64 ;
LAYER METAL3 ;
RECT 453.465 0.0 454.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[14]

PIN QA[14]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 463.285 496.265 464.355 496.905 ;
LAYER METAL2 ;
RECT 463.285 496.265 464.355 496.905 ;
LAYER METAL3 ;
RECT 463.285 496.265 464.355 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[14]

PIN DB[15]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 476.705 0.0 477.775 0.64 ;
LAYER METAL2 ;
RECT 476.705 0.0 477.775 0.64 ;
LAYER METAL3 ;
RECT 476.705 0.0 477.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[15]

PIN QA[15]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 486.525 496.265 487.595 496.905 ;
LAYER METAL2 ;
RECT 486.525 496.265 487.595 496.905 ;
LAYER METAL3 ;
RECT 486.525 496.265 487.595 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[15]

PIN DB[16]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 499.945 0.0 501.015 0.64 ;
LAYER METAL2 ;
RECT 499.945 0.0 501.015 0.64 ;
LAYER METAL3 ;
RECT 499.945 0.0 501.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[16]

PIN QA[16]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 509.765 496.265 510.835 496.905 ;
LAYER METAL2 ;
RECT 509.765 496.265 510.835 496.905 ;
LAYER METAL3 ;
RECT 509.765 496.265 510.835 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[16]

PIN DB[17]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 523.185 0.0 524.255 0.64 ;
LAYER METAL2 ;
RECT 523.185 0.0 524.255 0.64 ;
LAYER METAL3 ;
RECT 523.185 0.0 524.255 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[17]

PIN QA[17]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 533.005 496.265 534.075 496.905 ;
LAYER METAL2 ;
RECT 533.005 496.265 534.075 496.905 ;
LAYER METAL3 ;
RECT 533.005 496.265 534.075 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[17]

PIN DB[18]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 546.425 0.0 547.495 0.64 ;
LAYER METAL2 ;
RECT 546.425 0.0 547.495 0.64 ;
LAYER METAL3 ;
RECT 546.425 0.0 547.495 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[18]

PIN QA[18]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 556.245 496.265 557.315 496.905 ;
LAYER METAL2 ;
RECT 556.245 496.265 557.315 496.905 ;
LAYER METAL3 ;
RECT 556.245 496.265 557.315 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[18]

PIN DB[19]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 569.665 0.0 570.735 0.64 ;
LAYER METAL2 ;
RECT 569.665 0.0 570.735 0.64 ;
LAYER METAL3 ;
RECT 569.665 0.0 570.735 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[19]

PIN QA[19]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 579.485 496.265 580.555 496.905 ;
LAYER METAL2 ;
RECT 579.485 496.265 580.555 496.905 ;
LAYER METAL3 ;
RECT 579.485 496.265 580.555 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[19]

PIN DB[20]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 592.905 0.0 593.975 0.64 ;
LAYER METAL2 ;
RECT 592.905 0.0 593.975 0.64 ;
LAYER METAL3 ;
RECT 592.905 0.0 593.975 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[20]

PIN QA[20]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 602.725 496.265 603.795 496.905 ;
LAYER METAL2 ;
RECT 602.725 496.265 603.795 496.905 ;
LAYER METAL3 ;
RECT 602.725 496.265 603.795 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[20]

PIN DB[21]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 616.145 0.0 617.215 0.64 ;
LAYER METAL2 ;
RECT 616.145 0.0 617.215 0.64 ;
LAYER METAL3 ;
RECT 616.145 0.0 617.215 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[21]

PIN QA[21]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 625.965 496.265 627.035 496.905 ;
LAYER METAL2 ;
RECT 625.965 496.265 627.035 496.905 ;
LAYER METAL3 ;
RECT 625.965 496.265 627.035 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[21]

PIN DB[22]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 639.385 0.0 640.455 0.64 ;
LAYER METAL2 ;
RECT 639.385 0.0 640.455 0.64 ;
LAYER METAL3 ;
RECT 639.385 0.0 640.455 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[22]

PIN QA[22]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 649.205 496.265 650.275 496.905 ;
LAYER METAL2 ;
RECT 649.205 496.265 650.275 496.905 ;
LAYER METAL3 ;
RECT 649.205 496.265 650.275 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[22]

PIN DB[23]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 662.625 0.0 663.695 0.64 ;
LAYER METAL2 ;
RECT 662.625 0.0 663.695 0.64 ;
LAYER METAL3 ;
RECT 662.625 0.0 663.695 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[23]

PIN QA[23]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 672.445 496.265 673.515 496.905 ;
LAYER METAL2 ;
RECT 672.445 496.265 673.515 496.905 ;
LAYER METAL3 ;
RECT 672.445 496.265 673.515 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[23]

PIN VSS
DIRECTION INOUT ;
USE GROUND ;
PORT
LAYER METAL4 ;
RECT 279.475 0.0 283.475 496.905 ;
LAYER METAL4 ;
RECT 290.475 0.0 294.475 496.905 ;
LAYER METAL4 ;
RECT 301.475 0.0 305.475 496.905 ;
LAYER METAL4 ;
RECT 312.475 0.0 316.475 496.905 ;
LAYER METAL4 ;
RECT 323.475 0.0 327.475 496.905 ;
LAYER METAL4 ;
RECT 334.475 0.0 338.475 496.905 ;
LAYER METAL4 ;
RECT 343.945 0.0 347.945 496.905 ;
LAYER METAL4 ;
RECT 354.945 0.0 358.945 496.905 ;
LAYER METAL4 ;
RECT 365.945 0.0 369.945 496.905 ;
LAYER METAL4 ;
RECT 376.945 0.0 380.945 496.905 ;
LAYER METAL4 ;
RECT 387.945 0.0 391.945 496.905 ;
LAYER METAL4 ;
RECT 398.945 0.0 402.945 496.905 ;
LAYER METAL4 ;
RECT 267.855 0.0 271.855 496.905 ;
LAYER METAL4 ;
RECT 256.235 0.0 260.235 496.905 ;
LAYER METAL4 ;
RECT 244.615 0.0 248.615 496.905 ;
LAYER METAL4 ;
RECT 232.995 0.0 236.995 496.905 ;
LAYER METAL4 ;
RECT 221.375 0.0 225.375 496.905 ;
LAYER METAL4 ;
RECT 209.755 0.0 213.755 496.905 ;
LAYER METAL4 ;
RECT 198.135 0.0 202.135 496.905 ;
LAYER METAL4 ;
RECT 186.515 0.0 190.515 496.905 ;
LAYER METAL4 ;
RECT 174.895 0.0 178.895 496.905 ;
LAYER METAL4 ;
RECT 163.275 0.0 167.275 496.905 ;
LAYER METAL4 ;
RECT 151.655 0.0 155.655 496.905 ;
LAYER METAL4 ;
RECT 140.035 0.0 144.035 496.905 ;
LAYER METAL4 ;
RECT 128.415 0.0 132.415 496.905 ;
LAYER METAL4 ;
RECT 116.795 0.0 120.795 496.905 ;
LAYER METAL4 ;
RECT 105.175 0.0 109.175 496.905 ;
LAYER METAL4 ;
RECT 93.555 0.0 97.555 496.905 ;
LAYER METAL4 ;
RECT 81.935 0.0 85.935 496.905 ;
LAYER METAL4 ;
RECT 70.315 0.0 74.315 496.905 ;
LAYER METAL4 ;
RECT 58.695 0.0 62.695 496.905 ;
LAYER METAL4 ;
RECT 47.075 0.0 51.075 496.905 ;
LAYER METAL4 ;
RECT 35.455 0.0 39.455 496.905 ;
LAYER METAL4 ;
RECT 23.835 0.0 27.835 496.905 ;
LAYER METAL4 ;
RECT 12.215 0.0 16.215 496.905 ;
LAYER METAL4 ;
RECT 0.595 0.0 4.595 496.905 ;
LAYER METAL4 ;
RECT 410.565 0.0 414.565 496.905 ;
LAYER METAL4 ;
RECT 422.185 0.0 426.185 496.905 ;
LAYER METAL4 ;
RECT 433.805 0.0 437.805 496.905 ;
LAYER METAL4 ;
RECT 445.425 0.0 449.425 496.905 ;
LAYER METAL4 ;
RECT 457.045 0.0 461.045 496.905 ;
LAYER METAL4 ;
RECT 468.665 0.0 472.665 496.905 ;
LAYER METAL4 ;
RECT 480.285 0.0 484.285 496.905 ;
LAYER METAL4 ;
RECT 491.905 0.0 495.905 496.905 ;
LAYER METAL4 ;
RECT 503.525 0.0 507.525 496.905 ;
LAYER METAL4 ;
RECT 515.145 0.0 519.145 496.905 ;
LAYER METAL4 ;
RECT 526.765 0.0 530.765 496.905 ;
LAYER METAL4 ;
RECT 538.385 0.0 542.385 496.905 ;
LAYER METAL4 ;
RECT 550.005 0.0 554.005 496.905 ;
LAYER METAL4 ;
RECT 561.625 0.0 565.625 496.905 ;
LAYER METAL4 ;
RECT 573.245 0.0 577.245 496.905 ;
LAYER METAL4 ;
RECT 584.865 0.0 588.865 496.905 ;
LAYER METAL4 ;
RECT 596.485 0.0 600.485 496.905 ;
LAYER METAL4 ;
RECT 608.105 0.0 612.105 496.905 ;
LAYER METAL4 ;
RECT 619.725 0.0 623.725 496.905 ;
LAYER METAL4 ;
RECT 631.345 0.0 635.345 496.905 ;
LAYER METAL4 ;
RECT 642.965 0.0 646.965 496.905 ;
LAYER METAL4 ;
RECT 654.585 0.0 658.585 496.905 ;
LAYER METAL4 ;
RECT 666.205 0.0 670.205 496.905 ;
LAYER METAL4 ;
RECT 677.825 0.0 681.825 496.905 ;
END
END VSS

PIN VDD
DIRECTION INOUT ;
USE POWER ;
PORT
LAYER METAL4 ;
RECT 284.975 0.0 288.975 496.905 ;
LAYER METAL4 ;
RECT 295.975 0.0 299.975 496.905 ;
LAYER METAL4 ;
RECT 306.975 0.0 310.975 496.905 ;
LAYER METAL4 ;
RECT 317.975 0.0 321.975 496.905 ;
LAYER METAL4 ;
RECT 328.975 0.0 332.975 496.905 ;
LAYER METAL4 ;
RECT 349.445 0.0 353.445 496.905 ;
LAYER METAL4 ;
RECT 360.445 0.0 364.445 496.905 ;
LAYER METAL4 ;
RECT 371.445 0.0 375.445 496.905 ;
LAYER METAL4 ;
RECT 382.445 0.0 386.445 496.905 ;
LAYER METAL4 ;
RECT 393.445 0.0 397.445 496.905 ;
LAYER METAL4 ;
RECT 273.665 0.0 277.665 496.905 ;
LAYER METAL4 ;
RECT 262.045 0.0 266.045 496.905 ;
LAYER METAL4 ;
RECT 250.425 0.0 254.425 496.905 ;
LAYER METAL4 ;
RECT 238.805 0.0 242.805 496.905 ;
LAYER METAL4 ;
RECT 227.185 0.0 231.185 496.905 ;
LAYER METAL4 ;
RECT 215.565 0.0 219.565 496.905 ;
LAYER METAL4 ;
RECT 203.945 0.0 207.945 496.905 ;
LAYER METAL4 ;
RECT 192.325 0.0 196.325 496.905 ;
LAYER METAL4 ;
RECT 180.705 0.0 184.705 496.905 ;
LAYER METAL4 ;
RECT 169.085 0.0 173.085 496.905 ;
LAYER METAL4 ;
RECT 157.465 0.0 161.465 496.905 ;
LAYER METAL4 ;
RECT 145.845 0.0 149.845 496.905 ;
LAYER METAL4 ;
RECT 134.225 0.0 138.225 496.905 ;
LAYER METAL4 ;
RECT 122.605 0.0 126.605 496.905 ;
LAYER METAL4 ;
RECT 110.985 0.0 114.985 496.905 ;
LAYER METAL4 ;
RECT 99.365 0.0 103.365 496.905 ;
LAYER METAL4 ;
RECT 87.745 0.0 91.745 496.905 ;
LAYER METAL4 ;
RECT 76.125 0.0 80.125 496.905 ;
LAYER METAL4 ;
RECT 64.505 0.0 68.505 496.905 ;
LAYER METAL4 ;
RECT 52.885 0.0 56.885 496.905 ;
LAYER METAL4 ;
RECT 41.265 0.0 45.265 496.905 ;
LAYER METAL4 ;
RECT 29.645 0.0 33.645 496.905 ;
LAYER METAL4 ;
RECT 18.025 0.0 22.025 496.905 ;
LAYER METAL4 ;
RECT 6.405 0.0 10.405 496.905 ;
LAYER METAL4 ;
RECT 404.755 0.0 408.755 496.905 ;
LAYER METAL4 ;
RECT 416.375 0.0 420.375 496.905 ;
LAYER METAL4 ;
RECT 427.995 0.0 431.995 496.905 ;
LAYER METAL4 ;
RECT 439.615 0.0 443.615 496.905 ;
LAYER METAL4 ;
RECT 451.235 0.0 455.235 496.905 ;
LAYER METAL4 ;
RECT 462.855 0.0 466.855 496.905 ;
LAYER METAL4 ;
RECT 474.475 0.0 478.475 496.905 ;
LAYER METAL4 ;
RECT 486.095 0.0 490.095 496.905 ;
LAYER METAL4 ;
RECT 497.715 0.0 501.715 496.905 ;
LAYER METAL4 ;
RECT 509.335 0.0 513.335 496.905 ;
LAYER METAL4 ;
RECT 520.955 0.0 524.955 496.905 ;
LAYER METAL4 ;
RECT 532.575 0.0 536.575 496.905 ;
LAYER METAL4 ;
RECT 544.195 0.0 548.195 496.905 ;
LAYER METAL4 ;
RECT 555.815 0.0 559.815 496.905 ;
LAYER METAL4 ;
RECT 567.435 0.0 571.435 496.905 ;
LAYER METAL4 ;
RECT 579.055 0.0 583.055 496.905 ;
LAYER METAL4 ;
RECT 590.675 0.0 594.675 496.905 ;
LAYER METAL4 ;
RECT 602.295 0.0 606.295 496.905 ;
LAYER METAL4 ;
RECT 613.915 0.0 617.915 496.905 ;
LAYER METAL4 ;
RECT 625.535 0.0 629.535 496.905 ;
LAYER METAL4 ;
RECT 637.155 0.0 641.155 496.905 ;
LAYER METAL4 ;
RECT 648.775 0.0 652.775 496.905 ;
LAYER METAL4 ;
RECT 660.395 0.0 664.395 496.905 ;
LAYER METAL4 ;
RECT 672.015 0.0 676.015 496.905 ;
END
END VDD

OBS
LAYER VIA12 ;
RECT  0.000 0.000 682.420 496.905 ;
LAYER VIA23 ;
RECT  0.000 0.000 682.420 496.905 ;
LAYER VIA34 ;
RECT  0.000 0.000 682.420 496.905 ;
LAYER METAL1 ;
POLYGON 0.000 0.000 18.495 0.000 18.495 0.870 20.025 0.870 20.025 0.000
 41.735 0.000 41.735 0.870 43.265 0.870 43.265 0.000 64.975 0.000
 64.975 0.870 66.505 0.870 66.505 0.000 88.215 0.000 88.215 0.870
 89.745 0.870 89.745 0.000 111.455 0.000 111.455 0.870 112.985 0.870
 112.985 0.000 134.695 0.000 134.695 0.870 136.225 0.870 136.225 0.000
 157.935 0.000 157.935 0.870 159.465 0.870 159.465 0.000 181.175 0.000
 181.175 0.870 182.705 0.870 182.705 0.000 204.415 0.000 204.415 0.870
 205.945 0.870 205.945 0.000 227.655 0.000 227.655 0.870 229.185 0.870
 229.185 0.000 250.895 0.000 250.895 0.870 252.425 0.870 252.425 0.000
 274.135 0.000 274.135 0.870 275.665 0.870 275.665 0.000 296.875 0.000
 296.875 1.300 297.835 1.300 297.835 0.000 306.490 0.000 306.490 1.300
 307.450 1.300 307.450 0.000 323.220 0.000 323.220 0.870 325.245 0.870
 325.245 0.000 328.980 0.000 328.980 0.870 331.005 0.870 331.005 0.000
 334.740 0.000 334.740 0.870 336.765 0.870 336.765 0.000 340.500 0.000
 340.500 0.870 342.525 0.870 342.525 0.000 346.260 0.000 346.260 0.870
 348.285 0.870 348.285 0.000 351.785 0.000 351.785 0.870 353.895 0.870
 353.895 0.000 359.725 0.000 359.725 0.870 361.835 0.870 361.835 0.000
 367.665 0.000 367.665 0.870 369.775 0.870 369.775 0.000 378.435 0.000
 378.435 0.870 380.145 0.870 380.145 0.000 383.285 0.000 383.285 0.870
 384.995 0.870 384.995 0.000 406.755 0.000 406.755 0.870 408.285 0.870
 408.285 0.000 429.995 0.000 429.995 0.870 431.525 0.870 431.525 0.000
 453.235 0.000 453.235 0.870 454.765 0.870 454.765 0.000 476.475 0.000
 476.475 0.870 478.005 0.870 478.005 0.000 499.715 0.000 499.715 0.870
 501.245 0.870 501.245 0.000 522.955 0.000 522.955 0.870 524.485 0.870
 524.485 0.000 546.195 0.000 546.195 0.870 547.725 0.870 547.725 0.000
 569.435 0.000 569.435 0.870 570.965 0.870 570.965 0.000 592.675 0.000
 592.675 0.870 594.205 0.870 594.205 0.000 615.915 0.000 615.915 0.870
 617.445 0.870 617.445 0.000 639.155 0.000 639.155 0.870 640.685 0.870
 640.685 0.000 662.395 0.000 662.395 0.870 663.925 0.870 663.925 0.000
 682.420 0.000 682.420 496.905 673.745 496.905 673.745 496.035 672.215 496.035 672.215 496.905
 650.505 496.905 650.505 496.035 648.975 496.035 648.975 496.905 627.265 496.905
 627.265 496.035 625.735 496.035 625.735 496.905 604.025 496.905 604.025 496.035
 602.495 496.035 602.495 496.905 580.785 496.905 580.785 496.035 579.255 496.035
 579.255 496.905 557.545 496.905 557.545 496.035 556.015 496.035 556.015 496.905
 534.305 496.905 534.305 496.035 532.775 496.035 532.775 496.905 511.065 496.905
 511.065 496.035 509.535 496.035 509.535 496.905 487.825 496.905 487.825 496.035
 486.295 496.035 486.295 496.905 464.585 496.905 464.585 496.035 463.055 496.035
 463.055 496.905 441.345 496.905 441.345 496.035 439.815 496.035 439.815 496.905
 418.105 496.905 418.105 496.035 416.575 496.035 416.575 496.905 387.180 496.905
 387.180 495.605 386.220 495.605 386.220 496.905 377.775 496.905 377.775 495.605
 376.815 495.605 376.815 496.905 359.200 496.905 359.200 496.035 357.175 496.035
 357.175 496.905 353.440 496.905 353.440 496.035 351.415 496.035 351.415 496.905
 347.680 496.905 347.680 496.035 345.655 496.035 345.655 496.905 341.920 496.905
 341.920 496.035 339.895 496.035 339.895 496.905 336.160 496.905 336.160 496.035
 334.135 496.035 334.135 496.905 330.635 496.905 330.635 496.035 328.525 496.035
 328.525 496.905 322.695 496.905 322.695 496.035 320.585 496.035 320.585 496.905
 314.755 496.905 314.755 496.035 312.645 496.035 312.645 496.905 303.985 496.905
 303.985 496.035 302.275 496.035 302.275 496.905 299.135 496.905 299.135 496.035
 297.425 496.035 297.425 496.905 265.845 496.905 265.845 496.035 264.315 496.035
 264.315 496.905 242.605 496.905 242.605 496.035 241.075 496.035 241.075 496.905
 219.365 496.905 219.365 496.035 217.835 496.035 217.835 496.905 196.125 496.905
 196.125 496.035 194.595 496.035 194.595 496.905 172.885 496.905 172.885 496.035
 171.355 496.035 171.355 496.905 149.645 496.905 149.645 496.035 148.115 496.035
 148.115 496.905 126.405 496.905 126.405 496.035 124.875 496.035 124.875 496.905
 103.165 496.905 103.165 496.035 101.635 496.035 101.635 496.905 79.925 496.905
 79.925 496.035 78.395 496.035 78.395 496.905 56.685 496.905 56.685 496.035
 55.155 496.035 55.155 496.905 33.445 496.905 33.445 496.035 31.915 496.035
 31.915 496.905 10.205 496.905 10.205 496.035 8.675 496.035 8.675 496.905
 0.000 496.905 ;
LAYER METAL2 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 335.005 0.000 335.005 0.920 336.815 0.920 336.815 0.000 340.765 0.000
 340.765 0.920 342.575 0.920 342.575 0.000 346.525 0.000 346.525 0.920
 348.335 0.920 348.335 0.000 352.135 0.000 352.135 0.920 353.945 0.920
 353.945 0.000 360.075 0.000 360.075 0.920 361.885 0.920 361.885 0.000
 368.015 0.000 368.015 0.920 369.825 0.920 369.825 0.000 378.385 0.000
 378.385 0.920 380.195 0.920 380.195 0.000 383.235 0.000 383.235 0.920
 385.045 0.920 385.045 0.000 406.705 0.000 406.705 0.920 408.335 0.920
 408.335 0.000 429.945 0.000 429.945 0.920 431.575 0.920 431.575 0.000
 453.185 0.000 453.185 0.920 454.815 0.920 454.815 0.000 476.425 0.000
 476.425 0.920 478.055 0.920 478.055 0.000 499.665 0.000 499.665 0.920
 501.295 0.920 501.295 0.000 522.905 0.000 522.905 0.920 524.535 0.920
 524.535 0.000 546.145 0.000 546.145 0.920 547.775 0.920 547.775 0.000
 569.385 0.000 569.385 0.920 571.015 0.920 571.015 0.000 592.625 0.000
 592.625 0.920 594.255 0.920 594.255 0.000 615.865 0.000 615.865 0.920
 617.495 0.920 617.495 0.000 639.105 0.000 639.105 0.920 640.735 0.920
 640.735 0.000 662.345 0.000 662.345 0.920 663.975 0.920 663.975 0.000
 682.420 0.000 682.420 496.905 673.795 496.905 673.795 495.985 672.165 495.985 672.165 496.905
 650.555 496.905 650.555 495.985 648.925 495.985 648.925 496.905 627.315 496.905
 627.315 495.985 625.685 495.985 625.685 496.905 604.075 496.905 604.075 495.985
 602.445 495.985 602.445 496.905 580.835 496.905 580.835 495.985 579.205 495.985
 579.205 496.905 557.595 496.905 557.595 495.985 555.965 495.985 555.965 496.905
 534.355 496.905 534.355 495.985 532.725 495.985 532.725 496.905 511.115 496.905
 511.115 495.985 509.485 495.985 509.485 496.905 487.875 496.905 487.875 495.985
 486.245 495.985 486.245 496.905 464.635 496.905 464.635 495.985 463.005 495.985
 463.005 496.905 441.395 496.905 441.395 495.985 439.765 495.985 439.765 496.905
 418.155 496.905 418.155 495.985 416.525 495.985 416.525 496.905 387.230 496.905
 387.230 495.555 386.170 495.555 386.170 496.905 377.825 496.905 377.825 495.555
 376.765 495.555 376.765 496.905 358.935 496.905 358.935 495.985 357.125 495.985
 357.125 496.905 353.175 496.905 353.175 495.985 351.365 495.985 351.365 496.905
 347.415 496.905 347.415 495.985 345.605 495.985 345.605 496.905 341.655 496.905
 341.655 495.985 339.845 495.985 339.845 496.905 335.895 496.905 335.895 495.985
 334.085 495.985 334.085 496.905 330.285 496.905 330.285 495.985 328.475 495.985
 328.475 496.905 322.345 496.905 322.345 495.985 320.535 495.985 320.535 496.905
 314.405 496.905 314.405 495.985 312.595 495.985 312.595 496.905 304.035 496.905
 304.035 495.985 302.225 495.985 302.225 496.905 299.185 496.905 299.185 495.985
 297.375 495.985 297.375 496.905 265.895 496.905 265.895 495.985 264.265 495.985
 264.265 496.905 242.655 496.905 242.655 495.985 241.025 495.985 241.025 496.905
 219.415 496.905 219.415 495.985 217.785 495.985 217.785 496.905 196.175 496.905
 196.175 495.985 194.545 495.985 194.545 496.905 172.935 496.905 172.935 495.985
 171.305 495.985 171.305 496.905 149.695 496.905 149.695 495.985 148.065 495.985
 148.065 496.905 126.455 496.905 126.455 495.985 124.825 495.985 124.825 496.905
 103.215 496.905 103.215 495.985 101.585 495.985 101.585 496.905 79.975 496.905
 79.975 495.985 78.345 495.985 78.345 496.905 56.735 496.905 56.735 495.985
 55.105 495.985 55.105 496.905 33.495 496.905 33.495 495.985 31.865 495.985
 31.865 496.905 10.255 496.905 10.255 495.985 8.625 495.985 8.625 496.905
 0.000 496.905 ;
LAYER METAL3 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 335.005 0.000 335.005 0.920 336.815 0.920 336.815 0.000 340.765 0.000
 340.765 0.920 342.575 0.920 342.575 0.000 346.525 0.000 346.525 0.920
 348.335 0.920 348.335 0.000 352.135 0.000 352.135 0.920 353.945 0.920
 353.945 0.000 360.075 0.000 360.075 0.920 361.885 0.920 361.885 0.000
 368.015 0.000 368.015 0.920 369.825 0.920 369.825 0.000 378.385 0.000
 378.385 0.920 380.195 0.920 380.195 0.000 383.235 0.000 383.235 0.920
 385.045 0.920 385.045 0.000 406.705 0.000 406.705 0.920 408.335 0.920
 408.335 0.000 429.945 0.000 429.945 0.920 431.575 0.920 431.575 0.000
 453.185 0.000 453.185 0.920 454.815 0.920 454.815 0.000 476.425 0.000
 476.425 0.920 478.055 0.920 478.055 0.000 499.665 0.000 499.665 0.920
 501.295 0.920 501.295 0.000 522.905 0.000 522.905 0.920 524.535 0.920
 524.535 0.000 546.145 0.000 546.145 0.920 547.775 0.920 547.775 0.000
 569.385 0.000 569.385 0.920 571.015 0.920 571.015 0.000 592.625 0.000
 592.625 0.920 594.255 0.920 594.255 0.000 615.865 0.000 615.865 0.920
 617.495 0.920 617.495 0.000 639.105 0.000 639.105 0.920 640.735 0.920
 640.735 0.000 662.345 0.000 662.345 0.920 663.975 0.920 663.975 0.000
 682.420 0.000 682.420 496.905 673.795 496.905 673.795 495.985 672.165 495.985 672.165 496.905
 650.555 496.905 650.555 495.985 648.925 495.985 648.925 496.905 627.315 496.905
 627.315 495.985 625.685 495.985 625.685 496.905 604.075 496.905 604.075 495.985
 602.445 495.985 602.445 496.905 580.835 496.905 580.835 495.985 579.205 495.985
 579.205 496.905 557.595 496.905 557.595 495.985 555.965 495.985 555.965 496.905
 534.355 496.905 534.355 495.985 532.725 495.985 532.725 496.905 511.115 496.905
 511.115 495.985 509.485 495.985 509.485 496.905 487.875 496.905 487.875 495.985
 486.245 495.985 486.245 496.905 464.635 496.905 464.635 495.985 463.005 495.985
 463.005 496.905 441.395 496.905 441.395 495.985 439.765 495.985 439.765 496.905
 418.155 496.905 418.155 495.985 416.525 495.985 416.525 496.905 387.230 496.905
 387.230 495.555 386.170 495.555 386.170 496.905 377.825 496.905 377.825 495.555
 376.765 495.555 376.765 496.905 358.935 496.905 358.935 495.985 357.125 495.985
 357.125 496.905 353.175 496.905 353.175 495.985 351.365 495.985 351.365 496.905
 347.415 496.905 347.415 495.985 345.605 495.985 345.605 496.905 341.655 496.905
 341.655 495.985 339.845 495.985 339.845 496.905 335.895 496.905 335.895 495.985
 334.085 495.985 334.085 496.905 330.285 496.905 330.285 495.985 328.475 495.985
 328.475 496.905 322.345 496.905 322.345 495.985 320.535 495.985 320.535 496.905
 314.405 496.905 314.405 495.985 312.595 495.985 312.595 496.905 304.035 496.905
 304.035 495.985 302.225 495.985 302.225 496.905 299.185 496.905 299.185 495.985
 297.375 495.985 297.375 496.905 265.895 496.905 265.895 495.985 264.265 495.985
 264.265 496.905 242.655 496.905 242.655 495.985 241.025 495.985 241.025 496.905
 219.415 496.905 219.415 495.985 217.785 495.985 217.785 496.905 196.175 496.905
 196.175 495.985 194.545 495.985 194.545 496.905 172.935 496.905 172.935 495.985
 171.305 495.985 171.305 496.905 149.695 496.905 149.695 495.985 148.065 495.985
 148.065 496.905 126.455 496.905 126.455 495.985 124.825 495.985 124.825 496.905
 103.215 496.905 103.215 495.985 101.585 495.985 101.585 496.905 79.975 496.905
 79.975 495.985 78.345 495.985 78.345 496.905 56.735 496.905 56.735 495.985
 55.105 495.985 55.105 496.905 33.495 496.905 33.495 495.985 31.865 495.985
 31.865 496.905 10.255 496.905 10.255 495.985 8.625 495.985 8.625 496.905
 0.000 496.905 ;
END
END RAM1024
END LIBRARY
