************************************************************************
* auCdl Netlist:
*
* Library Name:  SMIC_MEMORY
* Top Cell Name: RAM256
* Version:  V0.2
* View Name:     schematic
* Netlisted on:  Mon Oct 31 21:44:15 CST 2022
************************************************************************
*.BIPOLAR
*.RESI = 2000
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM


************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELLDBL
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELLDBL BB VDD VSS
MM4 BB VSS VSS VSS N18 W=220.00N L=225.00N M=1
MM1 VSS VSS VSS VSS N18 W=705.00N L=180.00N M=1
MM7 VSS VSS VSS VSS N18 W=220.00N L=225.00N M=1
MM6 VDD VDD VDD VDD P18 W=220.000N L=200.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL_EDGE64
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL_EDGE64 DBL VDD VSS
XI0 DBL VDD VSS RAM256_BITCELLDBL
XI1 DBL VDD VSS RAM256_BITCELLDBL
XI2 DBL VDD VSS RAM256_BITCELLDBL
XI3 DBL VDD VSS RAM256_BITCELLDBL
XI4 DBL VDD VSS RAM256_BITCELLDBL
XI5 DBL VDD VSS RAM256_BITCELLDBL
XI6 DBL VDD VSS RAM256_BITCELLDBL
XI7 DBL VDD VSS RAM256_BITCELLDBL
XI8 DBL VDD VSS RAM256_BITCELLDBL
XI9 DBL VDD VSS RAM256_BITCELLDBL
XI10 DBL VDD VSS RAM256_BITCELLDBL
XI11 DBL VDD VSS RAM256_BITCELLDBL
XI12 DBL VDD VSS RAM256_BITCELLDBL
XI13 DBL VDD VSS RAM256_BITCELLDBL
XI14 DBL VDD VSS RAM256_BITCELLDBL
XI15 DBL VDD VSS RAM256_BITCELLDBL
XI16 DBL VDD VSS RAM256_BITCELLDBL
XI17 DBL VDD VSS RAM256_BITCELLDBL
XI18 DBL VDD VSS RAM256_BITCELLDBL
XI19 DBL VDD VSS RAM256_BITCELLDBL
XI20 DBL VDD VSS RAM256_BITCELLDBL
XI21 DBL VDD VSS RAM256_BITCELLDBL
XI22 DBL VDD VSS RAM256_BITCELLDBL
XI23 DBL VDD VSS RAM256_BITCELLDBL
XI24 DBL VDD VSS RAM256_BITCELLDBL
XI25 DBL VDD VSS RAM256_BITCELLDBL
XI26 DBL VDD VSS RAM256_BITCELLDBL
XI27 DBL VDD VSS RAM256_BITCELLDBL
XI28 DBL VDD VSS RAM256_BITCELLDBL
XI29 DBL VDD VSS RAM256_BITCELLDBL
XI30 DBL VDD VSS RAM256_BITCELLDBL
XI31 DBL VDD VSS RAM256_BITCELLDBL
XI32 DBL VDD VSS RAM256_BITCELLDBL
XI33 DBL VDD VSS RAM256_BITCELLDBL
XI34 DBL VDD VSS RAM256_BITCELLDBL
XI35 DBL VDD VSS RAM256_BITCELLDBL
XI36 DBL VDD VSS RAM256_BITCELLDBL
XI37 DBL VDD VSS RAM256_BITCELLDBL
XI38 DBL VDD VSS RAM256_BITCELLDBL
XI39 DBL VDD VSS RAM256_BITCELLDBL
XI40 DBL VDD VSS RAM256_BITCELLDBL
XI41 DBL VDD VSS RAM256_BITCELLDBL
XI42 DBL VDD VSS RAM256_BITCELLDBL
XI43 DBL VDD VSS RAM256_BITCELLDBL
XI44 DBL VDD VSS RAM256_BITCELLDBL
XI45 DBL VDD VSS RAM256_BITCELLDBL
XI46 DBL VDD VSS RAM256_BITCELLDBL
XI47 DBL VDD VSS RAM256_BITCELLDBL
XI48 DBL VDD VSS RAM256_BITCELLDBL
XI49 DBL VDD VSS RAM256_BITCELLDBL
XI50 DBL VDD VSS RAM256_BITCELLDBL
XI51 DBL VDD VSS RAM256_BITCELLDBL
XI52 DBL VDD VSS RAM256_BITCELLDBL
XI53 DBL VDD VSS RAM256_BITCELLDBL
XI54 DBL VDD VSS RAM256_BITCELLDBL
XI55 DBL VDD VSS RAM256_BITCELLDBL
XI56 DBL VDD VSS RAM256_BITCELLDBL
XI57 DBL VDD VSS RAM256_BITCELLDBL
XI58 DBL VDD VSS RAM256_BITCELLDBL
XI59 DBL VDD VSS RAM256_BITCELLDBL
XI60 DBL VDD VSS RAM256_BITCELLDBL
XI61 DBL VDD VSS RAM256_BITCELLDBL
XI62 DBL VDD VSS RAM256_BITCELLDBL
XI63 DBL VDD VSS RAM256_BITCELLDBL
XI64 NET12 VDD VSS RAM256_BITCELLDBL
XI65 NET12 VDD VSS RAM256_BITCELLDBL
XI66 NET18 VDD VSS RAM256_BITCELLDBL
XI67 DBL VDD VSS RAM256_BITCELLDBL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELLDUM
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELLDUM VSS WLA
MM4 VSS WLA VSS VSS N18 W=220.00N L=225.00N M=1
MM1 VSS VSS VSS VSS N18 W=705.00N L=180.00N M=1
MM7 VSS WLA VSS VSS N18 W=220.00N L=225.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_PCAP_DUMMY64
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_PCAP_DUMMY64 STWL[3] STWL[2] STWL[1] STWL[0] VSS WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 VSS WL[63] RAM256_BITCELLDUM
XI1 VSS WL[62] RAM256_BITCELLDUM
XI2 VSS WL[61] RAM256_BITCELLDUM
XI3 VSS WL[60] RAM256_BITCELLDUM
XI4 VSS WL[59] RAM256_BITCELLDUM
XI5 VSS WL[58] RAM256_BITCELLDUM
XI6 VSS WL[57] RAM256_BITCELLDUM
XI7 VSS WL[56] RAM256_BITCELLDUM
XI8 VSS WL[55] RAM256_BITCELLDUM
XI9 VSS WL[54] RAM256_BITCELLDUM
XI10 VSS WL[53] RAM256_BITCELLDUM
XI11 VSS WL[52] RAM256_BITCELLDUM
XI12 VSS WL[51] RAM256_BITCELLDUM
XI13 VSS WL[50] RAM256_BITCELLDUM
XI14 VSS WL[49] RAM256_BITCELLDUM
XI15 VSS WL[48] RAM256_BITCELLDUM
XI16 VSS WL[47] RAM256_BITCELLDUM
XI17 VSS WL[46] RAM256_BITCELLDUM
XI18 VSS WL[45] RAM256_BITCELLDUM
XI19 VSS WL[44] RAM256_BITCELLDUM
XI20 VSS WL[43] RAM256_BITCELLDUM
XI21 VSS WL[42] RAM256_BITCELLDUM
XI22 VSS WL[41] RAM256_BITCELLDUM
XI23 VSS WL[40] RAM256_BITCELLDUM
XI24 VSS WL[39] RAM256_BITCELLDUM
XI25 VSS WL[38] RAM256_BITCELLDUM
XI26 VSS WL[37] RAM256_BITCELLDUM
XI27 VSS WL[36] RAM256_BITCELLDUM
XI28 VSS WL[35] RAM256_BITCELLDUM
XI29 VSS WL[34] RAM256_BITCELLDUM
XI30 VSS WL[33] RAM256_BITCELLDUM
XI31 VSS WL[32] RAM256_BITCELLDUM
XI32 VSS WL[31] RAM256_BITCELLDUM
XI33 VSS WL[30] RAM256_BITCELLDUM
XI34 VSS WL[29] RAM256_BITCELLDUM
XI35 VSS WL[28] RAM256_BITCELLDUM
XI36 VSS WL[27] RAM256_BITCELLDUM
XI37 VSS WL[26] RAM256_BITCELLDUM
XI38 VSS WL[25] RAM256_BITCELLDUM
XI39 VSS WL[24] RAM256_BITCELLDUM
XI40 VSS WL[23] RAM256_BITCELLDUM
XI41 VSS WL[22] RAM256_BITCELLDUM
XI42 VSS WL[21] RAM256_BITCELLDUM
XI43 VSS WL[20] RAM256_BITCELLDUM
XI44 VSS WL[19] RAM256_BITCELLDUM
XI45 VSS WL[18] RAM256_BITCELLDUM
XI46 VSS WL[17] RAM256_BITCELLDUM
XI47 VSS WL[16] RAM256_BITCELLDUM
XI48 VSS WL[15] RAM256_BITCELLDUM
XI49 VSS WL[14] RAM256_BITCELLDUM
XI50 VSS WL[13] RAM256_BITCELLDUM
XI51 VSS WL[12] RAM256_BITCELLDUM
XI52 VSS WL[11] RAM256_BITCELLDUM
XI53 VSS WL[10] RAM256_BITCELLDUM
XI54 VSS WL[9] RAM256_BITCELLDUM
XI55 VSS WL[8] RAM256_BITCELLDUM
XI56 VSS WL[7] RAM256_BITCELLDUM
XI57 VSS WL[6] RAM256_BITCELLDUM
XI58 VSS WL[5] RAM256_BITCELLDUM
XI59 VSS WL[4] RAM256_BITCELLDUM
XI60 VSS WL[3] RAM256_BITCELLDUM
XI61 VSS STWL[3] RAM256_BITCELLDUM
XI62 VSS WL[2] RAM256_BITCELLDUM
XI63 VSS STWL[2] RAM256_BITCELLDUM
XI64 VSS WL[1] RAM256_BITCELLDUM
XI65 VSS STWL[1] RAM256_BITCELLDUM
XI66 VSS WL[0] RAM256_BITCELLDUM
XI67 VSS STWL[0] RAM256_BITCELLDUM
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_YMX4W_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_YMX4W_FLT BLW[3] BLW[2] BLW[1] BLW[0] BLXW[3] BLXW[2] BLXW[1] BLXW[0] CTRCLKW CTRCLKWX
+DATA VDD VSS YXW[3] YXW[2] YXW[1] YXW[0]
M0 VDD YXW[3] 7 VDD P18 L=1.8E-07 W=8E-07
M1 BLW[3] 7 VDD VDD P18 L=1.8E-07 W=1.5E-06
M2 9 YXW[2] VDD VDD P18 L=1.8E-07 W=8E-07
M3 BLXW[3] 7 BLW[3] VDD P18 L=1.8E-07 W=1.5E-06
M4 VDD 7 BLXW[3] VDD P18 L=1.8E-07 W=1.5E-06
M5 44 4 VDD VDD P18 L=1.8E-07 W=2.2E-07
M6 BLW[3] 7 VDD VDD P18 L=1.8E-07 W=1.5E-06
M7 8 CTRCLKWX 44 VDD P18 L=1.8E-07 W=2.2E-07
M8 BLXW[3] 7 BLW[3] VDD P18 L=1.8E-07 W=1.5E-06
M9 VDD 7 BLXW[3] VDD P18 L=1.8E-07 W=1.5E-06
M10 15 10 VDD VDD P18 L=1.8E-07 W=1.2E-06
M11 BLXW[2] 9 VDD VDD P18 L=1.8E-07 W=1.5E-06
M12 4 8 VDD VDD P18 L=1.8E-07 W=1.17E-06
M13 BLW[2] 9 BLXW[2] VDD P18 L=1.8E-07 W=1.5E-06
M14 VDD 8 4 VDD P18 L=1.8E-07 W=1.17E-06
M15 VDD 9 BLW[2] VDD P18 L=1.8E-07 W=1.5E-06
M16 VDD 11 10 VDD P18 L=5E-07 W=4E-07
M17 4 8 VDD VDD P18 L=1.8E-07 W=1.17E-06
M18 BLXW[2] 9 VDD VDD P18 L=1.8E-07 W=1.5E-06
M19 11 VSS VDD VDD P18 L=1.8E-07 W=4E-07
M20 8 CTRCLKW 32 VDD P18 L=1.8E-07 W=1E-06
M21 BLW[2] 9 BLXW[2] VDD P18 L=1.8E-07 W=1.5E-06
M22 32 CTRCLKW 8 VDD P18 L=1.8E-07 W=1E-06
M23 VDD 9 BLW[2] VDD P18 L=1.8E-07 W=1.5E-06
M24 VDD 13 14 VDD P18 L=1.8E-07 W=8E-07
M25 32 14 VDD VDD P18 L=1.8E-07 W=1.2E-06
M26 VDD 15 32 VDD P18 L=1.8E-07 W=1.2E-06
M27 34 15 VDD VDD P18 L=1.8E-07 W=1.2E-06
M28 16 CTRCLKW 34 VDD P18 L=1.8E-07 W=1E-06
M29 BLW[1] 20 VDD VDD P18 L=1.8E-07 W=1.5E-06
M30 VDD 13 34 VDD P18 L=1.8E-07 W=1.2E-06
M31 34 CTRCLKW 16 VDD P18 L=1.8E-07 W=1E-06
M32 BLXW[1] 20 BLW[1] VDD P18 L=1.8E-07 W=1.5E-06
M33 13 17 VDD VDD P18 L=1.8E-07 W=1.2E-06
M34 VDD 20 BLXW[1] VDD P18 L=1.8E-07 W=1.5E-06
M35 VDD 16 1 VDD P18 L=1.8E-07 W=1.17E-06
M36 BLW[1] 20 VDD VDD P18 L=1.8E-07 W=1.5E-06
M37 VDD 18 17 VDD P18 L=5E-07 W=4E-07
M38 1 16 VDD VDD P18 L=1.8E-07 W=1.17E-06
M39 BLXW[1] 20 BLW[1] VDD P18 L=1.8E-07 W=1.5E-06
M40 VDD DATA 18 VDD P18 L=1.8E-07 W=4E-07
M41 VDD 16 1 VDD P18 L=1.8E-07 W=1.17E-06
M42 VDD 20 BLXW[1] VDD P18 L=1.8E-07 W=1.5E-06
M43 BLXW[0] 21 VDD VDD P18 L=1.8E-07 W=1.5E-06
M44 45 CTRCLKWX 16 VDD P18 L=1.8E-07 W=2.2E-07
M45 BLW[0] 21 BLXW[0] VDD P18 L=1.8E-07 W=1.5E-06
M46 VDD 21 BLW[0] VDD P18 L=1.8E-07 W=1.5E-06
M47 VDD 1 45 VDD P18 L=1.8E-07 W=2.2E-07
M48 BLXW[0] 21 VDD VDD P18 L=1.8E-07 W=1.5E-06
M49 BLW[0] 21 BLXW[0] VDD P18 L=1.8E-07 W=1.5E-06
M50 VDD YXW[1] 20 VDD P18 L=1.8E-07 W=8E-07
M51 VDD 21 BLW[0] VDD P18 L=1.8E-07 W=1.5E-06
M52 21 YXW[0] VDD VDD P18 L=1.8E-07 W=8E-07
M53 BLW[3] 1 26 VSS N18 L=1.8E-07 W=1.75E-06
M54 VSS YXW[3] 7 VSS N18 L=1.8E-07 W=8E-07
M55 26 1 BLW[3] VSS N18 L=1.8E-07 W=1.75E-06
M56 9 YXW[2] VSS VSS N18 L=1.8E-07 W=8E-07
M57 VSS 7 26 VSS N18 L=1.8E-07 W=1.75E-06
M58 26 7 VSS VSS N18 L=1.8E-07 W=1.75E-06
M59 40 4 VSS VSS N18 L=1.8E-07 W=2.2E-07
M60 BLXW[3] 4 26 VSS N18 L=1.8E-07 W=1.75E-06
M61 8 CTRCLKW 40 VSS N18 L=1.8E-07 W=2.2E-07
M62 26 4 BLXW[3] VSS N18 L=1.8E-07 W=1.75E-06
M63 15 10 VSS VSS N18 L=1.8E-07 W=1.2E-06
M64 4 8 VSS VSS N18 L=1.8E-07 W=1.17E-06
M65 BLXW[2] 4 29 VSS N18 L=1.8E-07 W=1.75E-06
M66 VSS 8 4 VSS N18 L=1.8E-07 W=1.17E-06
M67 29 4 BLXW[2] VSS N18 L=1.8E-07 W=1.75E-06
M68 VSS 11 10 VSS N18 L=5E-07 W=4E-07
M69 4 8 VSS VSS N18 L=1.8E-07 W=1.17E-06
M70 VSS 9 29 VSS N18 L=1.8E-07 W=1.75E-06
M71 11 VSS VSS VSS N18 L=1.8E-07 W=4E-07
M72 29 9 VSS VSS N18 L=1.8E-07 W=1.75E-06
M73 8 CTRCLKWX 32 VSS N18 L=1.8E-07 W=1E-06
M74 BLW[2] 1 29 VSS N18 L=1.8E-07 W=1.75E-06
M75 32 CTRCLKWX 8 VSS N18 L=1.8E-07 W=1E-06
M76 29 1 BLW[2] VSS N18 L=1.8E-07 W=1.75E-06
M77 VSS 13 14 VSS N18 L=1.8E-07 W=8E-07
M78 41 14 VSS VSS N18 L=1.8E-07 W=1.2E-06
M79 32 15 41 VSS N18 L=1.8E-07 W=1.2E-06
M80 BLW[1] 1 33 VSS N18 L=1.8E-07 W=1.75E-06
M81 42 15 34 VSS N18 L=1.8E-07 W=1.2E-06
M82 16 CTRCLKWX 34 VSS N18 L=1.8E-07 W=1E-06
M83 33 1 BLW[1] VSS N18 L=1.8E-07 W=1.75E-06
M84 VSS 13 42 VSS N18 L=1.8E-07 W=1.2E-06
M85 34 CTRCLKWX 16 VSS N18 L=1.8E-07 W=1E-06
M86 VSS 20 33 VSS N18 L=1.8E-07 W=1.75E-06
M87 13 17 VSS VSS N18 L=1.8E-07 W=1.2E-06
M88 33 20 VSS VSS N18 L=1.8E-07 W=1.75E-06
M89 VSS 16 1 VSS N18 L=1.8E-07 W=1.17E-06
M90 BLXW[1] 4 33 VSS N18 L=1.8E-07 W=1.75E-06
M91 VSS 18 17 VSS N18 L=5E-07 W=4E-07
M92 1 16 VSS VSS N18 L=1.8E-07 W=1.17E-06
M93 33 4 BLXW[1] VSS N18 L=1.8E-07 W=1.75E-06
M94 VSS DATA 18 VSS N18 L=1.8E-07 W=4E-07
M95 VSS 16 1 VSS N18 L=1.8E-07 W=1.17E-06
M96 BLXW[0] 4 37 VSS N18 L=1.8E-07 W=1.75E-06
M97 43 CTRCLKW 16 VSS N18 L=1.8E-07 W=2.2E-07
M98 37 4 BLXW[0] VSS N18 L=1.8E-07 W=1.75E-06
M99 VSS 1 43 VSS N18 L=1.8E-07 W=2.2E-07
M100 VSS 21 37 VSS N18 L=1.8E-07 W=1.75E-06
M101 37 21 VSS VSS N18 L=1.8E-07 W=1.75E-06
M102 VSS YXW[1] 20 VSS N18 L=1.8E-07 W=8E-07
M103 BLW[0] 1 37 VSS N18 L=1.8E-07 W=1.75E-06
M104 21 YXW[0] VSS VSS N18 L=1.8E-07 W=8E-07
M105 37 1 BLW[0] VSS N18 L=1.8E-07 W=1.75E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_YMX4R_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_YMX4R_FLT BL[3] BL[2] BL[1] BL[0] BLX[3] BLX[2] BLX[1] BLX[0] DOUT VDD
+VSS YXR[3] YXR[2] YXR[1] YXR[0] CK1 CK4
M0 BL[0] 2 31 VDD P18 L=1.8E-07 W=5E-07
M1 VDD 2 1 VDD P18 L=1.8E-07 W=6.7E-07
M2 31 2 BL[0] VDD P18 L=1.8E-07 W=5E-07
M3 BL[0] 1 VDD VDD P18 L=1.8E-07 W=1E-06
M4 1 2 VDD VDD P18 L=1.8E-07 W=6.7E-07
M5 BL[0] 2 31 VDD P18 L=1.8E-07 W=5E-07
M6 BLX[0] 1 BL[0] VDD P18 L=1.8E-07 W=1E-06
M7 VDD 2 1 VDD P18 L=1.8E-07 W=6.7E-07
M8 VDD 1 BLX[0] VDD P18 L=1.8E-07 W=1E-06
M9 2 3 VDD VDD P18 L=1.8E-07 W=7E-07
M10 34 2 BLX[0] VDD P18 L=1.8E-07 W=5E-07
M11 BL[0] 1 VDD VDD P18 L=1.8E-07 W=1E-06
M12 VDD 3 2 VDD P18 L=1.8E-07 W=7E-07
M13 BLX[0] 2 34 VDD P18 L=1.8E-07 W=5E-07
M14 BLX[0] 1 BL[0] VDD P18 L=1.8E-07 W=1E-06
M15 34 2 BLX[0] VDD P18 L=1.8E-07 W=5E-07
M16 3 YXR[0] VDD VDD P18 L=1.8E-07 W=4E-07
M17 VDD 1 BLX[0] VDD P18 L=1.8E-07 W=1E-06
M18 BLX[1] 13 VDD VDD P18 L=1.8E-07 W=1E-06
M19 VDD YXR[1] 7 VDD P18 L=1.8E-07 W=4E-07
M20 BLX[1] 9 34 VDD P18 L=1.8E-07 W=5E-07
M21 31 11 8 VDD P18 L=1.8E-07 W=1.4E-06
M22 BL[1] 13 BLX[1] VDD P18 L=1.8E-07 W=1E-06
M23 VDD 8 10 VDD P18 L=2E-07 W=5.35E-07
M24 31 5 VDD VDD P18 L=1.8E-07 W=1E-06
M25 34 9 BLX[1] VDD P18 L=1.8E-07 W=5E-07
M26 9 7 VDD VDD P18 L=1.8E-07 W=7E-07
M27 8 11 31 VDD P18 L=1.8E-07 W=1.4E-06
M28 VDD 13 BL[1] VDD P18 L=1.8E-07 W=1E-06
M29 10 8 VDD VDD P18 L=2E-07 W=5.35E-07
M30 34 5 31 VDD P18 L=1.8E-07 W=1E-06
M31 BLX[1] 9 34 VDD P18 L=1.8E-07 W=5E-07
M32 VDD 7 9 VDD P18 L=1.8E-07 W=7E-07
M33 31 11 8 VDD P18 L=1.8E-07 W=1.4E-06
M34 BLX[1] 13 VDD VDD P18 L=1.8E-07 W=1E-06
M35 VDD 8 10 VDD P18 L=2E-07 W=5.35E-07
M36 VDD 5 34 VDD P18 L=1.8E-07 W=1E-06
M37 13 9 VDD VDD P18 L=1.8E-07 W=6.7E-07
M38 BL[1] 13 BLX[1] VDD P18 L=1.8E-07 W=1E-06
M39 8 10 VDD VDD P18 L=2E-07 W=5.35E-07
M40 31 5 VDD VDD P18 L=1.8E-07 W=1E-06
M41 31 9 BL[1] VDD P18 L=1.8E-07 W=5E-07
M42 VDD 9 13 VDD P18 L=1.8E-07 W=6.7E-07
M43 10 11 34 VDD P18 L=1.8E-07 W=1.4E-06
M44 VDD 13 BL[1] VDD P18 L=1.8E-07 W=1E-06
M45 34 5 31 VDD P18 L=1.8E-07 W=1E-06
M46 VDD 10 8 VDD P18 L=2E-07 W=5.35E-07
M47 BL[1] 9 31 VDD P18 L=1.8E-07 W=5E-07
M48 13 9 VDD VDD P18 L=1.8E-07 W=6.7E-07
M49 34 11 10 VDD P18 L=1.8E-07 W=1.4E-06
M50 VDD 5 34 VDD P18 L=1.8E-07 W=1E-06
M51 8 10 VDD VDD P18 L=2E-07 W=5.35E-07
M52 31 9 BL[1] VDD P18 L=1.8E-07 W=5E-07
M53 10 11 34 VDD P18 L=1.8E-07 W=1.4E-06
M54 17 CK4 VDD VDD P18 L=1.8E-07 W=4E-07
M55 VDD CK1 17 VDD P18 L=1.8E-07 W=4E-07
M56 BL[2] 21 31 VDD P18 L=1.8E-07 W=5E-07
M57 19 10 VDD VDD P18 L=1.8E-07 W=1.5E-06
M58 11 17 VDD VDD P18 L=1.8E-07 W=1.2E-06
M59 VDD 21 15 VDD P18 L=1.8E-07 W=6.7E-07
M60 31 21 BL[2] VDD P18 L=1.8E-07 W=5E-07
M61 BL[2] 15 VDD VDD P18 L=1.8E-07 W=1E-06
M62 VDD 18 19 VDD P18 L=1.8E-07 W=1.5E-06
M63 15 21 VDD VDD P18 L=1.8E-07 W=6.7E-07
M64 BL[2] 21 31 VDD P18 L=1.8E-07 W=5E-07
M65 BLX[2] 15 BL[2] VDD P18 L=1.8E-07 W=1E-06
M66 18 19 VDD VDD P18 L=1.8E-07 W=1.5E-06
M67 VDD 20 5 VDD P18 L=1.8E-07 W=1.6E-06
M68 VDD 21 15 VDD P18 L=1.8E-07 W=6.7E-07
M69 VDD 15 BLX[2] VDD P18 L=1.8E-07 W=1E-06
M70 VDD 8 18 VDD P18 L=1.8E-07 W=1.5E-06
M71 20 CK4 VDD VDD P18 L=1.8E-07 W=4E-07
M72 21 22 VDD VDD P18 L=1.8E-07 W=7E-07
M73 34 21 BLX[2] VDD P18 L=1.8E-07 W=5E-07
M74 BL[2] 15 VDD VDD P18 L=1.8E-07 W=1E-06
M75 VDD 22 21 VDD P18 L=1.8E-07 W=7E-07
M76 BLX[2] 21 34 VDD P18 L=1.8E-07 W=5E-07
M77 VDD CK1 23 VDD P18 L=1.8E-07 W=4E-07
M78 DOUT 18 VDD VDD P18 L=1.8E-07 W=2E-06
M79 BLX[2] 15 BL[2] VDD P18 L=1.8E-07 W=1E-06
M80 34 21 BLX[2] VDD P18 L=1.8E-07 W=5E-07
M81 22 YXR[2] VDD VDD P18 L=1.8E-07 W=4E-07
M82 12 23 VDD VDD P18 L=1.8E-07 W=1.2E-06
M83 VDD 18 DOUT VDD P18 L=1.8E-07 W=2E-06
M84 VDD 15 BLX[2] VDD P18 L=1.8E-07 W=1E-06
M85 BLX[3] 28 VDD VDD P18 L=1.8E-07 W=1E-06
M86 VDD YXR[3] 26 VDD P18 L=1.8E-07 W=4E-07
M87 BLX[3] 27 34 VDD P18 L=1.8E-07 W=5E-07
M88 BL[3] 28 BLX[3] VDD P18 L=1.8E-07 W=1E-06
M89 34 27 BLX[3] VDD P18 L=1.8E-07 W=5E-07
M90 27 26 VDD VDD P18 L=1.8E-07 W=7E-07
M91 VDD 28 BL[3] VDD P18 L=1.8E-07 W=1E-06
M92 BLX[3] 27 34 VDD P18 L=1.8E-07 W=5E-07
M93 VDD 26 27 VDD P18 L=1.8E-07 W=7E-07
M94 BLX[3] 28 VDD VDD P18 L=1.8E-07 W=1E-06
M95 28 27 VDD VDD P18 L=1.8E-07 W=6.7E-07
M96 BL[3] 28 BLX[3] VDD P18 L=1.8E-07 W=1E-06
M97 31 27 BL[3] VDD P18 L=1.8E-07 W=5E-07
M98 VDD 27 28 VDD P18 L=1.8E-07 W=6.7E-07
M99 VDD 28 BL[3] VDD P18 L=1.8E-07 W=1E-06
M100 BL[3] 27 31 VDD P18 L=1.8E-07 W=5E-07
M101 28 27 VDD VDD P18 L=1.8E-07 W=6.7E-07
M102 31 27 BL[3] VDD P18 L=1.8E-07 W=5E-07
M103 VSS 2 1 VSS N18 L=1.8E-07 W=6.7E-07
M104 1 2 VSS VSS N18 L=1.8E-07 W=6.7E-07
M105 VSS 2 1 VSS N18 L=1.8E-07 W=6.7E-07
M106 2 3 VSS VSS N18 L=1.8E-07 W=6E-07
M107 VSS 3 2 VSS N18 L=1.8E-07 W=6E-07
M108 3 YXR[0] VSS VSS N18 L=1.8E-07 W=4E-07
M109 VSS YXR[1] 7 VSS N18 L=1.8E-07 W=4E-07
M110 10 8 36 VSS N18 L=2E-07 W=3E-06
M111 43 5 VSS VSS N18 L=1.8E-07 W=2E-06
M112 36 12 43 VSS N18 L=1.8E-07 W=2E-06
M113 9 7 VSS VSS N18 L=1.8E-07 W=6E-07
M114 36 8 10 VSS N18 L=2E-07 W=3E-06
M115 VSS 7 9 VSS N18 L=1.8E-07 W=6E-07
M116 8 10 36 VSS N18 L=2E-07 W=3E-06
M117 13 9 VSS VSS N18 L=1.8E-07 W=6.7E-07
M118 36 10 8 VSS N18 L=2E-07 W=3E-06
M119 VSS 9 13 VSS N18 L=1.8E-07 W=6.7E-07
M120 13 9 VSS VSS N18 L=1.8E-07 W=6.7E-07
M121 44 CK4 17 VSS N18 L=1.8E-07 W=4E-07
M122 VSS CK1 44 VSS N18 L=1.8E-07 W=4E-07
M123 11 17 VSS VSS N18 L=1.8E-07 W=1.2E-06
M124 45 10 19 VSS N18 L=1.8E-07 W=1.5E-06
M125 VSS 21 15 VSS N18 L=1.8E-07 W=6.7E-07
M126 VSS 18 45 VSS N18 L=1.8E-07 W=1.5E-06
M127 15 21 VSS VSS N18 L=1.8E-07 W=6.7E-07
M128 46 19 VSS VSS N18 L=1.8E-07 W=1.5E-06
M129 VSS 20 5 VSS N18 L=1.8E-07 W=1.2E-06
M130 VSS 21 15 VSS N18 L=1.8E-07 W=6.7E-07
M131 18 8 46 VSS N18 L=1.8E-07 W=1.5E-06
M132 20 CK4 VSS VSS N18 L=1.8E-07 W=8E-07
M133 21 22 VSS VSS N18 L=1.8E-07 W=6E-07
M134 VSS CK1 23 VSS N18 L=1.8E-07 W=4E-07
M135 VSS 22 21 VSS N18 L=1.8E-07 W=6E-07
M136 DOUT 18 VSS VSS N18 L=1.8E-07 W=1E-06
M137 22 YXR[2] VSS VSS N18 L=1.8E-07 W=4E-07
M138 12 23 VSS VSS N18 L=1.8E-07 W=1.2E-06
M139 VSS 18 DOUT VSS N18 L=1.8E-07 W=1E-06
M140 VSS YXR[3] 26 VSS N18 L=1.8E-07 W=4E-07
M141 27 26 VSS VSS N18 L=1.8E-07 W=6E-07
M142 VSS 26 27 VSS N18 L=1.8E-07 W=6E-07
M143 28 27 VSS VSS N18 L=1.8E-07 W=6.7E-07
M144 VSS 27 28 VSS N18 L=1.8E-07 W=6.7E-07
M145 28 27 VSS VSS N18 L=1.8E-07 W=6.7E-07
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_YMX4SAWR_AB
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_YMX4SAWR_AB BLA[3] BLA[2] BLA[1] BLA[0] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[3] BLXA[2]
+BLXA[1] BLXA[0] BLXB[3] BLXB[2] BLXB[1] BLXB[0] CK1 CK4 CTRCLK CTRCLKX
+DATA QA VDD VSS YXR[3] YXR[2] YXR[1] YXR[0] YXW[3] YXW[2]
+YXW[1] YXW[0]
XYMUXW BLB[3] BLB[2] BLB[1] BLB[0] BLXB[3] BLXB[2] BLXB[1] BLXB[0] CTRCLK 
+ CTRCLKX DATA VDD VSS YXW[3] YXW[2] YXW[1] YXW[0] / RAM256_YMX4W_FLT
XYMUXR BLA[3] BLA[2] BLA[1] BLA[0] BLXA[3] BLXA[2] BLXA[1] BLXA[0] QA VDD VSS 
+ YXR[3] YXR[2] YXR[1] YXR[0] CK1 CK4 / RAM256_YMX4R_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL8T
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL8T BA BB BXA BXB VDD VSS WLA WLB
MM0 BCN BC VSS VSS N18 W=705.00N L=180.00N M=1
MM4 BB WLB BC VSS N18 W=220.00N L=225.00N M=1
MM1 BC BCN VSS VSS N18 W=705.00N L=180.00N M=1
MM2 BXA WLA BCN VSS N18 W=220.00N L=225.00N M=1
MM3 BA WLA BC VSS N18 W=220.00N L=225.00N M=1
MM7 BXB WLB BCN VSS N18 W=220.00N L=225.00N M=1
MM5 BCN BC VDD VDD P18 W=220.000N L=200.00N M=1
MM6 BC BCN VDD VDD P18 W=220.000N L=200.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL2X2
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL2X2 BA[1] BA[0] BB[1] BB[0] BXA[1] BXA[0] BXB[1] BXB[0] VDD VSS
+WLA[1] WLA[0] WLB[1] WLB[0]
XI8 BA[0] BB[0] BXA[0] BXB[0] VDD VSS WLA[0] WLB[0] RAM256_BITCELL8T
XI11 BA[1] BB[1] BXA[1] BXB[1] VDD VSS WLA[1] WLB[1] RAM256_BITCELL8T
XI9 BA[0] BB[0] BXA[0] BXB[0] VDD VSS WLA[1] WLB[1] RAM256_BITCELL8T
XI10 BA[1] BB[1] BXA[1] BXB[1] VDD VSS WLA[0] WLB[0] RAM256_BITCELL8T
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL32X2N
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL32X2N BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[31] WLA[30] WLB[31] WLB[30] RAM256_BITCELL2X2
XI1 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[29] WLA[28] WLB[29] WLB[28] RAM256_BITCELL2X2
XI2 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[27] WLA[26] WLB[27] WLB[26] RAM256_BITCELL2X2
XI3 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[25] WLA[24] WLB[25] WLB[24] RAM256_BITCELL2X2
XI4 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[23] WLA[22] WLB[23] WLB[22] RAM256_BITCELL2X2
XI5 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[21] WLA[20] WLB[21] WLB[20] RAM256_BITCELL2X2
XI6 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[19] WLA[18] WLB[19] WLB[18] RAM256_BITCELL2X2
XI7 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[17] WLA[16] WLB[17] WLB[16] RAM256_BITCELL2X2
XI8 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[15] WLA[14] WLB[15] WLB[14] RAM256_BITCELL2X2
XI9 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[13] WLA[12] WLB[13] WLB[12] RAM256_BITCELL2X2
XI10 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[11] WLA[10] WLB[11] WLB[10] RAM256_BITCELL2X2
XI11 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[9] WLA[8] WLB[9] WLB[8] RAM256_BITCELL2X2
XI12 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[7] WLA[6] WLB[7] WLB[6] RAM256_BITCELL2X2
XI13 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[5] WLA[4] WLB[5] WLB[4] RAM256_BITCELL2X2
XI14 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[3] WLA[2] WLB[3] WLB[2] RAM256_BITCELL2X2
XI15 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[1] WLA[0] WLB[1] WLB[0] RAM256_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL64X2
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL64X2 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL32X2N
XI1 BLXA[1] BLXA[0] BLXB[1] BLXB[0] BLA[1] BLA[0] BLB[1] BLB[0] VDD VSS
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] RAM256_BITCELL32X2N
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL2X2_STWL
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL2X2_STWL BA0 BXA0 VDD VSS WLA[3] WLA[2] WLA[1] WLA[0] WLB[3] WLB[2] WLB[1] WLB[0]
XI8 BA0 NET54 BXA0 NET53 VDD VSS WLA[0] WLB[0] RAM256_BITCELL8T
XI11 BA3 NET46 BXA3 NET45 VDD VSS WLA[3] WLB[3] RAM256_BITCELL8T
XI9 NET64 NET54 NET63 NET53 VDD VSS WLA[1] WLB[1] RAM256_BITCELL8T
XI10 NET64 NET46 NET63 NET45 VDD VSS WLA[2] WLB[2] RAM256_BITCELL8T
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL64X2ABR
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL64X2ABR BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] RDWLA[3] RDWLA[2]
+RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL64X2
XI1 BLA[1] BLXA[1] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RAM256_BITCELL2X2_STWL
XI2 BLA[0] BLXA[0] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RAM256_BITCELL2X2_STWL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_ARRAY_X64Y4D1
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_ARRAY_X64Y4D1 CLKB CLKXB DATAB DOUTA RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 BLA[3] BLA[2] BLA[1] BLA[0] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[3] BLXA[2]
+BLXA[1] BLXA[0] BLXB[3] BLXB[2] BLXB[1] BLXB[0] SACK1A SACK4A CLKB CLKXB
+DATAB DOUTA VDD VSS YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2]
+YXB[1] YXB[0] RAM256_YMX4SAWR_AB
XI1 BLA[3] BLA[2] BLB[3] BLB[2] BLXA[3] BLXA[2] BLXB[3] BLXB[2] VSS VSS
+VSS VSS RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL64X2ABR
XI2 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VSS VSS
+VSS VSS RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL64X2ABR
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_BITCELL64X2ABR_MID
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_BITCELL64X2ABR_MID BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] RDWLA[3] RDWLA[2]
+RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL64X2
XI1 BLA[1] BLXA[1] VDD VSS RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] RAM256_BITCELL2X2_STWL
XI2 BLA[0] BLXA[0] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RAM256_BITCELL2X2_STWL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_ARRAY_X64Y4D1_MD
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_ARRAY_X64Y4D1_MD CLKB CLKXB DATAB DOUTA RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2]
+RDWLB_MID[1] RDWLB_MID[0] SACK1A SACK4A VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2]
+YXB[1] YXB[0]
XI0 BLA[3] BLA[2] BLA[1] BLA[0] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[3] BLXA[2]
+BLXA[1] BLXA[0] BLXB[3] BLXB[2] BLXB[1] BLXB[0] SACK1A SACK4A CLKB CLKXB
+DATAB DOUTA VDD VSS YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2]
+YXB[1] YXB[0] RAM256_YMX4SAWR_AB
XI1 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VSS VSS
+VSS VSS RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL64X2ABR
XI2 BLA[3] BLA[2] BLB[3] BLB[2] BLXA[3] BLXA[2] BLXB[3] BLXB[2] VSS VSS
+VSS VSS VSS VSS VSS VSS RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] RAM256_BITCELL64X2ABR_MID
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_ARRAY_X64Y4D12_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_ARRAY_X64Y4D12_RIGHT CLKB CLKXB DATAB[11] DATAB[10] DATAB[9] DATAB[8] DATAB[7] DATAB[6] DATAB[5] DATAB[4]
+DATAB[3] DATAB[2] DATAB[1] DATAB[0] DBL DOUTA[11] DOUTA[10] DOUTA[9] DOUTA[8] DOUTA[7]
+DOUTA[6] DOUTA[5] DOUTA[4] DOUTA[3] DOUTA[2] DOUTA[1] DOUTA[0] SACK1A SACK4A STWLA
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 DBL VDD VSS RAM256_BITCELL_EDGE64
XI1 VSS VSS VSS VSS VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] RAM256_PCAP_DUMMY64
XI2 CLKB CLKXB DATAB[11] DOUTA[11] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI3 CLKB CLKXB DATAB[10] DOUTA[10] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI4 CLKB CLKXB DATAB[9] DOUTA[9] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI5 CLKB CLKXB DATAB[8] DOUTA[8] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI6 CLKB CLKXB DATAB[7] DOUTA[7] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI7 CLKB CLKXB DATAB[6] DOUTA[6] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI8 CLKB CLKXB DATAB[5] DOUTA[5] VSS STWLA STWLA VSS VSS STWLA
+STWLA VSS SACK1A SACK4A VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2]
+YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1_MD
XI9 CLKB CLKXB DATAB[4] DOUTA[4] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI10 CLKB CLKXB DATAB[3] DOUTA[3] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI11 CLKB CLKXB DATAB[2] DOUTA[2] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI12 CLKB CLKXB DATAB[1] DOUTA[1] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI13 CLKB CLKXB DATAB[0] DOUTA[0] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_ARRAY_X64Y4D12_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_ARRAY_X64Y4D12_LEFT CLKB CLKXB DATAB[11] DATAB[10] DATAB[9] DATAB[8] DATAB[7] DATAB[6] DATAB[5] DATAB[4]
+DATAB[3] DATAB[2] DATAB[1] DATAB[0] DBL DOUTA[11] DOUTA[10] DOUTA[9] DOUTA[8] DOUTA[7]
+DOUTA[6] DOUTA[5] DOUTA[4] DOUTA[3] DOUTA[2] DOUTA[1] DOUTA[0] SACK1A SACK4A STWLA
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 DBL VDD VSS RAM256_BITCELL_EDGE64
XI1 VSS VSS VSS VSS VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] RAM256_PCAP_DUMMY64
XI2 CLKB CLKXB DATAB[11] DOUTA[11] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI3 CLKB CLKXB DATAB[10] DOUTA[10] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI4 CLKB CLKXB DATAB[9] DOUTA[9] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI5 CLKB CLKXB DATAB[8] DOUTA[8] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI6 CLKB CLKXB DATAB[7] DOUTA[7] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI7 CLKB CLKXB DATAB[6] DOUTA[6] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI8 CLKB CLKXB DATAB[5] DOUTA[5] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI9 CLKB CLKXB DATAB[4] DOUTA[4] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI10 CLKB CLKXB DATAB[3] DOUTA[3] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI11 CLKB CLKXB DATAB[2] DOUTA[2] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI12 CLKB CLKXB DATAB[1] DOUTA[1] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
XI13 CLKB CLKXB DATAB[0] DOUTA[0] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXA[3] YXA[2] YXA[1] YXA[0] YXB[3] YXB[2] YXB[1] YXB[0] RAM256_ARRAY_X64Y4D1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_SOP_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_SOP_FLT DBLA EMCLKA S[1] S[0] STWLA VDD VSS
M0 8 EMCLKA VDD VDD P18 L=1.8E-07 W=1.6E-06
M1 VDD EMCLKA 8 VDD P18 L=1.8E-07 W=1.6E-06
M2 STWLA 8 VDD VDD P18 L=1.8E-07 W=2E-06
M3 VDD 8 STWLA VDD P18 L=1.8E-07 W=2E-06
M4 STWLA 8 VDD VDD P18 L=1.8E-07 W=2E-06
M5 VDD 8 STWLA VDD P18 L=1.8E-07 W=2E-06
M6 STWLA 8 VDD VDD P18 L=1.8E-07 W=2E-06
M7 VDD S[0] 11 VDD P18 L=1.8E-07 W=1.2E-06
M8 10 S[1] VDD VDD P18 L=1.8E-07 W=1.2E-06
M9 VDD 10 3 VDD P18 L=1.8E-07 W=1.2E-06
M10 4 10 VDD VDD P18 L=1.8E-07 W=1.2E-06
M11 VDD 11 4 VDD P18 L=1.8E-07 W=1.2E-06
M12 19 11 VDD VDD P18 L=1.8E-07 W=1.2E-06
M13 5 10 19 VDD P18 L=1.8E-07 W=1.2E-06
M14 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M15 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M16 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M17 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M18 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M19 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M20 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M21 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M22 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M23 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M24 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M25 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M26 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M27 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M28 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M29 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M30 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M31 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M32 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M33 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M34 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M35 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M36 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M37 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M38 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M39 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M40 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M41 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M42 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M43 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M44 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M45 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M46 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M47 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M48 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M49 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M50 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M51 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M52 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M53 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M54 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M55 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M56 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M57 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M58 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M59 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M60 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M61 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M62 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M63 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M64 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M65 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M66 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M67 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M68 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M69 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M70 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M71 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M72 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M73 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M74 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M75 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M76 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M77 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M78 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M79 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M80 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M81 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M82 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M83 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M84 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M85 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M86 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M87 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M88 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M89 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M90 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M91 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M92 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M93 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M94 VSS S[0] 11 VSS N18 L=1.8E-07 W=1.2E-06
M95 10 S[1] VSS VSS N18 L=1.8E-07 W=1.2E-06
M96 VSS 10 3 VSS N18 L=1.8E-07 W=1.2E-06
M97 18 10 VSS VSS N18 L=1.8E-07 W=1.2E-06
M98 4 11 18 VSS N18 L=1.8E-07 W=1.2E-06
M99 5 11 VSS VSS N18 L=1.8E-07 W=1.2E-06
M100 VSS 10 5 VSS N18 L=1.8E-07 W=1.2E-06
M101 STWLA 8 VSS VSS N18 L=1.8E-07 W=1E-06
M102 VSS 8 STWLA VSS N18 L=1.8E-07 W=1E-06
M103 STWLA 8 VSS VSS N18 L=1.8E-07 W=1E-06
M104 VSS 8 STWLA VSS N18 L=1.8E-07 W=1E-06
M105 STWLA 8 VSS VSS N18 L=1.8E-07 W=1E-06
M106 8 EMCLKA VSS VSS N18 L=1.8E-07 W=8E-07
M107 VSS EMCLKA 8 VSS N18 L=1.8E-07 W=8E-07
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_SOP_W_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_SOP_W_FLT DBLB EMCLKB S[1] S[0] VDD VSS
M0 VDD S[0] 9 VDD P18 L=1.8E-07 W=1.2E-06
M1 8 S[1] VDD VDD P18 L=1.8E-07 W=1.2E-06
M2 VDD 8 3 VDD P18 L=1.8E-07 W=1.2E-06
M3 4 8 VDD VDD P18 L=1.8E-07 W=1.2E-06
M4 VDD 9 4 VDD P18 L=1.8E-07 W=1.2E-06
M5 17 9 VDD VDD P18 L=1.8E-07 W=1.2E-06
M6 5 8 17 VDD P18 L=1.8E-07 W=1.2E-06
M7 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M8 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M9 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M10 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M11 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M12 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M13 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M14 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M15 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M16 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M17 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M18 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M19 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M20 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M21 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M22 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M23 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M24 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M25 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M26 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M27 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M28 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M29 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M30 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M31 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M32 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M33 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M34 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M35 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M36 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M37 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M38 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M39 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M40 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M41 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M42 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M43 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M44 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M45 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M46 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M47 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M48 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M49 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M50 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M51 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M52 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M53 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M54 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M55 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M56 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M57 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M58 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M59 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M60 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M61 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M62 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M63 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M64 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M65 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M66 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M67 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M68 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M69 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M70 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M71 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M72 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M73 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M74 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M75 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M76 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M77 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M78 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M79 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M80 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M81 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M82 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M83 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M84 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M85 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M86 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M87 VSS S[0] 9 VSS N18 L=1.8E-07 W=1.2E-06
M88 8 S[1] VSS VSS N18 L=1.8E-07 W=1.2E-06
M89 VSS 8 3 VSS N18 L=1.8E-07 W=1.2E-06
M90 16 8 VSS VSS N18 L=1.8E-07 W=1.2E-06
M91 4 9 16 VSS N18 L=1.8E-07 W=1.2E-06
M92 5 9 VSS VSS N18 L=1.8E-07 W=1.2E-06
M93 VSS 8 5 VSS N18 L=1.8E-07 W=1.2E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_LEAFCELL_PX4_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_LEAFCELL_PX4_FLT A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] VDD VSS
M0 19 2 VDD VDD P18 L=1.8E-07 W=1E-06
M1 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M2 3 CLK 19 VDD P18 L=1.8E-07 W=8.35E-07
M3 VDD 4 19 VDD P18 L=1.8E-07 W=1E-06
M4 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M5 19 CLK 3 VDD P18 L=1.8E-07 W=8.35E-07
M6 VDD PX[0] 3 VDD P18 L=1E-06 W=2.2E-07
M7 4 A[0] VDD VDD P18 L=1.8E-07 W=4E-07
M8 19 4 VDD VDD P18 L=1.8E-07 W=1E-06
M9 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M10 3 CLK 19 VDD P18 L=1.8E-07 W=8.35E-07
M11 VDD A[0] 4 VDD P18 L=1.8E-07 W=4E-07
M12 VDD 2 19 VDD P18 L=1.8E-07 W=1E-06
M13 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M14 20 2 VDD VDD P18 L=1.8E-07 W=1E-06
M15 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M16 9 4 VDD VDD P18 L=1.8E-07 W=4E-07
M17 10 PX[1] VDD VDD P18 L=1E-06 W=2.2E-07
M18 20 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M19 VDD 9 20 VDD P18 L=1.8E-07 W=1E-06
M20 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M21 VDD 4 9 VDD P18 L=1.8E-07 W=4E-07
M22 10 CLK 20 VDD P18 L=1.8E-07 W=8.35E-07
M23 20 9 VDD VDD P18 L=1.8E-07 W=1E-06
M24 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M25 20 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M26 VDD 2 20 VDD P18 L=1.8E-07 W=1E-06
M27 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M28 21 11 VDD VDD P18 L=1.8E-07 W=1E-06
M29 PX[2] 12 VDD VDD P18 L=1.8E-07 W=2.5E-06
M30 12 CLK 21 VDD P18 L=1.8E-07 W=8.35E-07
M31 VDD 4 21 VDD P18 L=1.8E-07 W=1E-06
M32 VDD 12 PX[2] VDD P18 L=1.8E-07 W=2.5E-06
M33 21 CLK 12 VDD P18 L=1.8E-07 W=8.35E-07
M34 VDD PX[2] 12 VDD P18 L=1E-06 W=2.2E-07
M35 2 A[1] VDD VDD P18 L=1.8E-07 W=4E-07
M36 21 4 VDD VDD P18 L=1.8E-07 W=1E-06
M37 PX[2] 12 VDD VDD P18 L=1.8E-07 W=2.5E-06
M38 12 CLK 21 VDD P18 L=1.8E-07 W=8.35E-07
M39 VDD A[1] 2 VDD P18 L=1.8E-07 W=4E-07
M40 VDD 11 21 VDD P18 L=1.8E-07 W=1E-06
M41 VDD 12 PX[2] VDD P18 L=1.8E-07 W=2.5E-06
M42 22 11 VDD VDD P18 L=1.8E-07 W=1E-06
M43 PX[3] 16 VDD VDD P18 L=1.8E-07 W=2.5E-06
M44 11 2 VDD VDD P18 L=1.8E-07 W=4E-07
M45 16 PX[3] VDD VDD P18 L=1E-06 W=2.2E-07
M46 22 CLK 16 VDD P18 L=1.8E-07 W=8.35E-07
M47 VDD 9 22 VDD P18 L=1.8E-07 W=1E-06
M48 VDD 16 PX[3] VDD P18 L=1.8E-07 W=2.5E-06
M49 VDD 2 11 VDD P18 L=1.8E-07 W=4E-07
M50 16 CLK 22 VDD P18 L=1.8E-07 W=8.35E-07
M51 22 9 VDD VDD P18 L=1.8E-07 W=1E-06
M52 PX[3] 16 VDD VDD P18 L=1.8E-07 W=2.5E-06
M53 22 CLK 16 VDD P18 L=1.8E-07 W=8.35E-07
M54 VDD 11 22 VDD P18 L=1.8E-07 W=1E-06
M55 VDD 16 PX[3] VDD P18 L=1.8E-07 W=2.5E-06
M56 23 2 VSS VSS N18 L=1.8E-07 W=1E-06
M57 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M58 19 4 23 VSS N18 L=1.8E-07 W=1E-06
M59 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M60 19 CLKX 3 VSS N18 L=1.8E-07 W=1.25E-06
M61 VSS PX[0] 3 VSS N18 L=1E-06 W=2.2E-07
M62 4 A[0] VSS VSS N18 L=1.8E-07 W=4E-07
M63 24 4 19 VSS N18 L=1.8E-07 W=1E-06
M64 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M65 3 CLKX 19 VSS N18 L=1.8E-07 W=1.25E-06
M66 VSS A[0] 4 VSS N18 L=1.8E-07 W=4E-07
M67 VSS 2 24 VSS N18 L=1.8E-07 W=1E-06
M68 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M69 25 2 VSS VSS N18 L=1.8E-07 W=1E-06
M70 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M71 9 4 VSS VSS N18 L=1.8E-07 W=4E-07
M72 10 PX[1] VSS VSS N18 L=1E-06 W=2.2E-07
M73 20 CLKX 10 VSS N18 L=1.8E-07 W=1.25E-06
M74 20 9 25 VSS N18 L=1.8E-07 W=1E-06
M75 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
M76 VSS 4 9 VSS N18 L=1.8E-07 W=4E-07
M77 10 CLKX 20 VSS N18 L=1.8E-07 W=1.25E-06
M78 26 9 20 VSS N18 L=1.8E-07 W=1E-06
M79 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M80 VSS 2 26 VSS N18 L=1.8E-07 W=1E-06
M81 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
M82 27 11 VSS VSS N18 L=1.8E-07 W=1E-06
M83 PX[2] 12 VSS VSS N18 L=1.8E-07 W=1E-06
M84 21 4 27 VSS N18 L=1.8E-07 W=1E-06
M85 VSS 12 PX[2] VSS N18 L=1.8E-07 W=1E-06
M86 21 CLKX 12 VSS N18 L=1.8E-07 W=1.25E-06
M87 VSS PX[2] 12 VSS N18 L=1E-06 W=2.2E-07
M88 2 A[1] VSS VSS N18 L=1.8E-07 W=4E-07
M89 28 4 21 VSS N18 L=1.8E-07 W=1E-06
M90 PX[2] 12 VSS VSS N18 L=1.8E-07 W=1E-06
M91 12 CLKX 21 VSS N18 L=1.8E-07 W=1.25E-06
M92 VSS A[1] 2 VSS N18 L=1.8E-07 W=4E-07
M93 VSS 11 28 VSS N18 L=1.8E-07 W=1E-06
M94 VSS 12 PX[2] VSS N18 L=1.8E-07 W=1E-06
M95 29 11 VSS VSS N18 L=1.8E-07 W=1E-06
M96 PX[3] 16 VSS VSS N18 L=1.8E-07 W=1E-06
M97 11 2 VSS VSS N18 L=1.8E-07 W=4E-07
M98 16 PX[3] VSS VSS N18 L=1E-06 W=2.2E-07
M99 22 CLKX 16 VSS N18 L=1.8E-07 W=1.25E-06
M100 22 9 29 VSS N18 L=1.8E-07 W=1E-06
M101 VSS 16 PX[3] VSS N18 L=1.8E-07 W=1E-06
M102 VSS 2 11 VSS N18 L=1.8E-07 W=4E-07
M103 16 CLKX 22 VSS N18 L=1.8E-07 W=1.25E-06
M104 30 9 22 VSS N18 L=1.8E-07 W=1E-06
M105 PX[3] 16 VSS VSS N18 L=1.8E-07 W=1E-06
M106 VSS 11 30 VSS N18 L=1.8E-07 W=1E-06
M107 VSS 16 PX[3] VSS N18 L=1.8E-07 W=1E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_LEAFCELL_PX2_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_LEAFCELL_PX2_FLT A[0] CLK CLKX PX[1] PX[0] VDD VSS
M0 12 2 VDD VDD P18 L=1.8E-07 W=1E-06
M1 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M2 3 CLK 12 VDD P18 L=1.8E-07 W=8.35E-07
M3 VDD VDD 12 VDD P18 L=1.8E-07 W=1E-06
M4 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M5 12 CLK 3 VDD P18 L=1.8E-07 W=8.35E-07
M6 VDD PX[0] 3 VDD P18 L=1E-06 W=2.2E-07
M7 2 A[0] VDD VDD P18 L=1.8E-07 W=4E-07
M8 12 VDD VDD VDD P18 L=1.8E-07 W=1E-06
M9 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M10 3 CLK 12 VDD P18 L=1.8E-07 W=8.35E-07
M11 VDD A[0] 2 VDD P18 L=1.8E-07 W=4E-07
M12 VDD 2 12 VDD P18 L=1.8E-07 W=1E-06
M13 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M14 13 8 VDD VDD P18 L=1.8E-07 W=1E-06
M15 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M16 8 2 VDD VDD P18 L=1.8E-07 W=4E-07
M17 10 PX[1] VDD VDD P18 L=1E-06 W=2.2E-07
M18 13 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M19 VDD VDD 13 VDD P18 L=1.8E-07 W=1E-06
M20 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M21 VDD 2 8 VDD P18 L=1.8E-07 W=4E-07
M22 10 CLK 13 VDD P18 L=1.8E-07 W=8.35E-07
M23 13 VDD VDD VDD P18 L=1.8E-07 W=1E-06
M24 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M25 13 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M26 VDD 8 13 VDD P18 L=1.8E-07 W=1E-06
M27 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M28 14 2 VSS VSS N18 L=1.8E-07 W=1E-06
M29 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M30 12 VDD 14 VSS N18 L=1.8E-07 W=1E-06
M31 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M32 12 CLKX 3 VSS N18 L=1.8E-07 W=1.25E-06
M33 VSS PX[0] 3 VSS N18 L=1E-06 W=2.2E-07
M34 2 A[0] VSS VSS N18 L=1.8E-07 W=4E-07
M35 15 VDD 12 VSS N18 L=1.8E-07 W=1E-06
M36 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M37 3 CLKX 12 VSS N18 L=1.8E-07 W=1.25E-06
M38 VSS A[0] 2 VSS N18 L=1.8E-07 W=4E-07
M39 VSS 2 15 VSS N18 L=1.8E-07 W=1E-06
M40 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M41 16 8 VSS VSS N18 L=1.8E-07 W=1E-06
M42 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M43 8 2 VSS VSS N18 L=1.8E-07 W=4E-07
M44 10 PX[1] VSS VSS N18 L=1E-06 W=2.2E-07
M45 13 CLKX 10 VSS N18 L=1.8E-07 W=1.25E-06
M46 13 VDD 16 VSS N18 L=1.8E-07 W=1E-06
M47 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
M48 VSS 2 8 VSS N18 L=1.8E-07 W=4E-07
M49 10 CLKX 13 VSS N18 L=1.8E-07 W=1.25E-06
M50 17 VDD 13 VSS N18 L=1.8E-07 W=1E-06
M51 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M52 VSS 8 17 VSS N18 L=1.8E-07 W=1E-06
M53 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_FPREDEC_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_FPREDEC_FLT A[0] A[1] A[2] CLK CLKX FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] VDD VSS WLCKX
M0 1 A[0] VDD VDD P18 L=1.8E-07 W=8E-07
M1 31 1 VDD VDD P18 L=1.8E-07 W=1E-06
M2 FCKX[2] 4 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M3 FCKX[2] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M4 4 CLK 31 VDD P18 L=1.8E-07 W=1.6E-06
M5 VDD 5 31 VDD P18 L=1.8E-07 W=1E-06
M6 WLCKX 4 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M7 VDD 6 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M8 VDD 6 4 VDD P18 L=1E-06 W=2.2E-07
M9 31 8 VDD VDD P18 L=1.8E-07 W=1E-06
M10 FCKX[2] 4 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M11 FCKX[2] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M12 VDD 4 6 VDD P18 L=1.8E-07 W=1.6E-06
M13 WLCKX 4 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M14 VDD 6 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M15 9 10 VDD VDD P18 L=1.8E-07 W=1.6E-06
M16 FCKX[3] 10 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M17 FCKX[3] 9 VDD VDD P18 L=1.8E-07 W=1.25E-06
M18 10 9 VDD VDD P18 L=1E-06 W=2.2E-07
M19 VDD 8 33 VDD P18 L=1.8E-07 W=1E-06
M20 WLCKX 10 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M21 VDD 9 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M22 33 5 VDD VDD P18 L=1.8E-07 W=1E-06
M23 FCKX[3] 10 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M24 FCKX[3] 9 VDD VDD P18 L=1.8E-07 W=1.25E-06
M25 33 CLK 10 VDD P18 L=1.8E-07 W=1.6E-06
M26 VDD 11 33 VDD P18 L=1.8E-07 W=1E-06
M27 WLCKX 10 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M28 VDD 9 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M29 35 11 VDD VDD P18 L=1.8E-07 W=1E-06
M30 FCKX[1] 12 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M31 FCKX[1] 13 VDD VDD P18 L=1.8E-07 W=1.25E-06
M32 11 1 VDD VDD P18 L=1.8E-07 W=8E-07
M33 12 CLK 35 VDD P18 L=1.8E-07 W=1.6E-06
M34 VDD 5 35 VDD P18 L=1.8E-07 W=1E-06
M35 WLCKX 12 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M36 VDD 13 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M37 VDD 13 12 VDD P18 L=1E-06 W=2.2E-07
M38 35 14 VDD VDD P18 L=1.8E-07 W=1E-06
M39 FCKX[1] 12 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M40 FCKX[1] 13 VDD VDD P18 L=1.8E-07 W=1.25E-06
M41 14 A[1] VDD VDD P18 L=1.8E-07 W=8E-07
M42 VDD 12 13 VDD P18 L=1.8E-07 W=1.6E-06
M43 WLCKX 12 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M44 VDD 13 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M45 15 17 VDD VDD P18 L=1.8E-07 W=1.6E-06
M46 FCKX[0] 17 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M47 FCKX[0] 15 VDD VDD P18 L=1.8E-07 W=1.25E-06
M48 17 15 VDD VDD P18 L=1E-06 W=2.2E-07
M49 VDD 14 37 VDD P18 L=1.8E-07 W=1E-06
M50 WLCKX 17 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M51 VDD 15 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M52 37 5 VDD VDD P18 L=1.8E-07 W=1E-06
M53 FCKX[0] 17 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M54 FCKX[0] 15 VDD VDD P18 L=1.8E-07 W=1.25E-06
M55 37 CLK 17 VDD P18 L=1.8E-07 W=1.6E-06
M56 VDD 1 37 VDD P18 L=1.8E-07 W=1E-06
M57 WLCKX 17 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M58 VDD 15 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M59 39 1 VDD VDD P18 L=1.8E-07 W=1E-06
M60 FCKX[4] 18 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M61 FCKX[4] 20 VDD VDD P18 L=1.8E-07 W=1.25E-06
M62 18 CLK 39 VDD P18 L=1.8E-07 W=1.6E-06
M63 VDD 19 39 VDD P18 L=1.8E-07 W=1E-06
M64 WLCKX 18 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M65 VDD 20 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M66 VDD 20 18 VDD P18 L=1E-06 W=2.2E-07
M67 39 14 VDD VDD P18 L=1.8E-07 W=1E-06
M68 FCKX[4] 18 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M69 FCKX[4] 20 VDD VDD P18 L=1.8E-07 W=1.25E-06
M70 VDD 18 20 VDD P18 L=1.8E-07 W=1.6E-06
M71 WLCKX 18 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M72 VDD 20 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M73 8 14 VDD VDD P18 L=1.8E-07 W=8E-07
M74 21 22 VDD VDD P18 L=1.8E-07 W=1.6E-06
M75 FCKX[5] 22 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M76 FCKX[5] 21 VDD VDD P18 L=1.8E-07 W=1.25E-06
M77 22 21 VDD VDD P18 L=1E-06 W=2.2E-07
M78 VDD 14 41 VDD P18 L=1.8E-07 W=1E-06
M79 WLCKX 22 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M80 VDD 21 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M81 5 A[2] VDD VDD P18 L=1.8E-07 W=8E-07
M82 41 19 VDD VDD P18 L=1.8E-07 W=1E-06
M83 FCKX[5] 22 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M84 FCKX[5] 21 VDD VDD P18 L=1.8E-07 W=1.25E-06
M85 41 CLK 22 VDD P18 L=1.8E-07 W=1.6E-06
M86 VDD 11 41 VDD P18 L=1.8E-07 W=1E-06
M87 WLCKX 22 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M88 VDD 21 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M89 43 11 VDD VDD P18 L=1.8E-07 W=1E-06
M90 FCKX[7] 24 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M91 FCKX[7] 25 VDD VDD P18 L=1.8E-07 W=1.25E-06
M92 24 CLK 43 VDD P18 L=1.8E-07 W=1.6E-06
M93 VDD 19 43 VDD P18 L=1.8E-07 W=1E-06
M94 WLCKX 24 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M95 VDD 25 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M96 VDD 25 24 VDD P18 L=1E-06 W=2.2E-07
M97 43 8 VDD VDD P18 L=1.8E-07 W=1E-06
M98 FCKX[7] 24 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M99 FCKX[7] 25 VDD VDD P18 L=1.8E-07 W=1.25E-06
M100 VDD 24 25 VDD P18 L=1.8E-07 W=1.6E-06
M101 WLCKX 24 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M102 VDD 25 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M103 26 27 VDD VDD P18 L=1.8E-07 W=1.6E-06
M104 FCKX[6] 27 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M105 FCKX[6] 26 VDD VDD P18 L=1.8E-07 W=1.25E-06
M106 27 26 VDD VDD P18 L=1E-06 W=2.2E-07
M107 VDD 8 45 VDD P18 L=1.8E-07 W=1E-06
M108 WLCKX 27 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M109 VDD 26 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M110 45 19 VDD VDD P18 L=1.8E-07 W=1E-06
M111 FCKX[6] 27 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M112 FCKX[6] 26 VDD VDD P18 L=1.8E-07 W=1.25E-06
M113 45 CLK 27 VDD P18 L=1.8E-07 W=1.6E-06
M114 19 5 VDD VDD P18 L=1.8E-07 W=8E-07
M115 VDD 1 45 VDD P18 L=1.8E-07 W=1E-06
M116 WLCKX 27 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M117 VDD 26 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M118 47 1 VSS VSS N18 L=1.8E-07 W=1E-06
M119 FCKX[2] 6 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M120 4 CLKX 31 VSS N18 L=1.8E-07 W=1.6E-06
M121 48 5 47 VSS N18 L=1.8E-07 W=1E-06
M122 WLCKX 6 FCKX[2] VSS N18 L=1.8E-07 W=1.25E-06
M123 VSS 6 4 VSS N18 L=1E-06 W=2.2E-07
M124 31 8 48 VSS N18 L=1.8E-07 W=1E-06
M125 FCKX[2] 6 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M126 1 A[0] VSS VSS N18 L=1.8E-07 W=8E-07
M127 VSS 4 6 VSS N18 L=1.8E-07 W=1.6E-06
M128 WLCKX 6 FCKX[2] VSS N18 L=1.8E-07 W=1.25E-06
M129 9 10 VSS VSS N18 L=1.8E-07 W=1.6E-06
M130 FCKX[3] 9 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M131 10 9 VSS VSS N18 L=1E-06 W=2.2E-07
M132 49 8 33 VSS N18 L=1.8E-07 W=1E-06
M133 WLCKX 9 FCKX[3] VSS N18 L=1.8E-07 W=1.25E-06
M134 11 1 VSS VSS N18 L=1.8E-07 W=8E-07
M135 50 5 49 VSS N18 L=1.8E-07 W=1E-06
M136 FCKX[3] 9 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M137 33 CLKX 10 VSS N18 L=1.8E-07 W=1.6E-06
M138 VSS 11 50 VSS N18 L=1.8E-07 W=1E-06
M139 WLCKX 9 FCKX[3] VSS N18 L=1.8E-07 W=1.25E-06
M140 51 11 VSS VSS N18 L=1.8E-07 W=1E-06
M141 FCKX[1] 13 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M142 12 CLKX 35 VSS N18 L=1.8E-07 W=1.6E-06
M143 52 5 51 VSS N18 L=1.8E-07 W=1E-06
M144 WLCKX 13 FCKX[1] VSS N18 L=1.8E-07 W=1.25E-06
M145 VSS 13 12 VSS N18 L=1E-06 W=2.2E-07
M146 35 14 52 VSS N18 L=1.8E-07 W=1E-06
M147 FCKX[1] 13 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M148 VSS 12 13 VSS N18 L=1.8E-07 W=1.6E-06
M149 WLCKX 13 FCKX[1] VSS N18 L=1.8E-07 W=1.25E-06
M150 15 17 VSS VSS N18 L=1.8E-07 W=1.6E-06
M151 FCKX[0] 15 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M152 17 15 VSS VSS N18 L=1E-06 W=2.2E-07
M153 53 14 37 VSS N18 L=1.8E-07 W=1E-06
M154 WLCKX 15 FCKX[0] VSS N18 L=1.8E-07 W=1.25E-06
M155 14 A[1] VSS VSS N18 L=1.8E-07 W=8E-07
M156 54 5 53 VSS N18 L=1.8E-07 W=1E-06
M157 FCKX[0] 15 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M158 37 CLKX 17 VSS N18 L=1.8E-07 W=1.6E-06
M159 VSS 1 54 VSS N18 L=1.8E-07 W=1E-06
M160 WLCKX 15 FCKX[0] VSS N18 L=1.8E-07 W=1.25E-06
M161 55 1 VSS VSS N18 L=1.8E-07 W=1E-06
M162 FCKX[4] 20 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M163 18 CLKX 39 VSS N18 L=1.8E-07 W=1.6E-06
M164 8 14 VSS VSS N18 L=1.8E-07 W=8E-07
M165 56 19 55 VSS N18 L=1.8E-07 W=1E-06
M166 WLCKX 20 FCKX[4] VSS N18 L=1.8E-07 W=1.25E-06
M167 VSS 20 18 VSS N18 L=1E-06 W=2.2E-07
M168 39 14 56 VSS N18 L=1.8E-07 W=1E-06
M169 FCKX[4] 20 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M170 VSS 18 20 VSS N18 L=1.8E-07 W=1.6E-06
M171 WLCKX 20 FCKX[4] VSS N18 L=1.8E-07 W=1.25E-06
M172 21 22 VSS VSS N18 L=1.8E-07 W=1.6E-06
M173 FCKX[5] 21 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M174 22 21 VSS VSS N18 L=1E-06 W=2.2E-07
M175 57 14 41 VSS N18 L=1.8E-07 W=1E-06
M176 WLCKX 21 FCKX[5] VSS N18 L=1.8E-07 W=1.25E-06
M177 58 19 57 VSS N18 L=1.8E-07 W=1E-06
M178 FCKX[5] 21 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M179 41 CLKX 22 VSS N18 L=1.8E-07 W=1.6E-06
M180 VSS 11 58 VSS N18 L=1.8E-07 W=1E-06
M181 WLCKX 21 FCKX[5] VSS N18 L=1.8E-07 W=1.25E-06
M182 59 11 VSS VSS N18 L=1.8E-07 W=1E-06
M183 FCKX[7] 25 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M184 5 A[2] VSS VSS N18 L=1.8E-07 W=8E-07
M185 24 CLKX 43 VSS N18 L=1.8E-07 W=1.6E-06
M186 60 19 59 VSS N18 L=1.8E-07 W=1E-06
M187 WLCKX 25 FCKX[7] VSS N18 L=1.8E-07 W=1.25E-06
M188 VSS 25 24 VSS N18 L=1E-06 W=2.2E-07
M189 43 8 60 VSS N18 L=1.8E-07 W=1E-06
M190 FCKX[7] 25 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M191 VSS 24 25 VSS N18 L=1.8E-07 W=1.6E-06
M192 WLCKX 25 FCKX[7] VSS N18 L=1.8E-07 W=1.25E-06
M193 19 5 VSS VSS N18 L=1.8E-07 W=8E-07
M194 26 27 VSS VSS N18 L=1.8E-07 W=1.6E-06
M195 FCKX[6] 26 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M196 27 26 VSS VSS N18 L=1E-06 W=2.2E-07
M197 61 8 45 VSS N18 L=1.8E-07 W=1E-06
M198 WLCKX 26 FCKX[6] VSS N18 L=1.8E-07 W=1.25E-06
M199 62 19 61 VSS N18 L=1.8E-07 W=1E-06
M200 FCKX[6] 26 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M201 45 CLKX 27 VSS N18 L=1.8E-07 W=1.6E-06
M202 VSS 1 62 VSS N18 L=1.8E-07 W=1E-06
M203 WLCKX 26 FCKX[6] VSS N18 L=1.8E-07 W=1.25E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_YPREDEC4_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_YPREDEC4_FLT A[0] A[1] CLK CLKX VDD VSS YCKX YX[3] YX[2] YX[1] YX[0]
M0 20 1 VDD VDD P18 L=1.8E-07 W=1E-06
M1 YX[0] 4 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M2 YX[0] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M3 4 CLK 20 VDD P18 L=1.8E-07 W=1.6E-06
M4 VDD 5 20 VDD P18 L=1.8E-07 W=1E-06
M5 YCKX 4 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M6 VDD 6 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M7 VDD 6 4 VDD P18 L=1E-06 W=2.2E-07
M8 YX[0] 4 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M9 YX[0] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M10 VDD A[0] 1 VDD P18 L=1.8E-07 W=8E-07
M11 VDD 4 6 VDD P18 L=1.8E-07 W=1.6E-06
M12 YCKX 4 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M13 VDD 6 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M14 10 1 VDD VDD P18 L=1.8E-07 W=8E-07
M15 8 9 VDD VDD P18 L=1.8E-07 W=1.6E-06
M16 YX[1] 9 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M17 YX[1] 8 VDD VDD P18 L=1.8E-07 W=1.25E-06
M18 9 8 VDD VDD P18 L=1E-06 W=2.2E-07
M19 YCKX 9 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M20 VDD 8 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M21 23 5 VDD VDD P18 L=1.8E-07 W=1E-06
M22 YX[1] 9 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M23 YX[1] 8 VDD VDD P18 L=1.8E-07 W=1.25E-06
M24 23 CLK 9 VDD P18 L=1.8E-07 W=1.6E-06
M25 VDD 10 23 VDD P18 L=1.8E-07 W=1E-06
M26 YCKX 9 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M27 VDD 8 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M28 24 10 VDD VDD P18 L=1.8E-07 W=1E-06
M29 YX[3] 11 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M30 YX[3] 13 VDD VDD P18 L=1.8E-07 W=1.25E-06
M31 11 CLK 24 VDD P18 L=1.8E-07 W=1.6E-06
M32 VDD 12 24 VDD P18 L=1.8E-07 W=1E-06
M33 YCKX 11 YX[3] VDD P18 L=1.8E-07 W=1.25E-06
M34 VDD 13 YX[3] VDD P18 L=1.8E-07 W=1.25E-06
M35 VDD 13 11 VDD P18 L=1E-06 W=2.2E-07
M36 YX[3] 11 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M37 YX[3] 13 VDD VDD P18 L=1.8E-07 W=1.25E-06
M38 VDD A[1] 5 VDD P18 L=1.8E-07 W=8E-07
M39 VDD 11 13 VDD P18 L=1.8E-07 W=1.6E-06
M40 YCKX 11 YX[3] VDD P18 L=1.8E-07 W=1.25E-06
M41 VDD 13 YX[3] VDD P18 L=1.8E-07 W=1.25E-06
M42 12 5 VDD VDD P18 L=1.8E-07 W=8E-07
M43 15 16 VDD VDD P18 L=1.8E-07 W=1.6E-06
M44 YX[2] 16 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M45 YX[2] 15 VDD VDD P18 L=1.8E-07 W=1.25E-06
M46 16 15 VDD VDD P18 L=1E-06 W=2.2E-07
M47 YCKX 16 YX[2] VDD P18 L=1.8E-07 W=1.25E-06
M48 VDD 15 YX[2] VDD P18 L=1.8E-07 W=1.25E-06
M49 27 12 VDD VDD P18 L=1.8E-07 W=1E-06
M50 YX[2] 16 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M51 YX[2] 15 VDD VDD P18 L=1.8E-07 W=1.25E-06
M52 27 CLK 16 VDD P18 L=1.8E-07 W=1.6E-06
M53 VDD 1 27 VDD P18 L=1.8E-07 W=1E-06
M54 YCKX 16 YX[2] VDD P18 L=1.8E-07 W=1.25E-06
M55 VDD 15 YX[2] VDD P18 L=1.8E-07 W=1.25E-06
M56 28 1 VSS VSS N18 L=1.8E-07 W=1E-06
M57 YX[0] 6 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M58 4 CLKX 20 VSS N18 L=1.8E-07 W=1.6E-06
M59 20 5 28 VSS N18 L=1.8E-07 W=1E-06
M60 YCKX 6 YX[0] VSS N18 L=1.8E-07 W=1.25E-06
M61 VSS 6 4 VSS N18 L=1E-06 W=2.2E-07
M62 YX[0] 6 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M63 VSS A[0] 1 VSS N18 L=1.8E-07 W=8E-07
M64 VSS 4 6 VSS N18 L=1.8E-07 W=1.6E-06
M65 YCKX 6 YX[0] VSS N18 L=1.8E-07 W=1.25E-06
M66 10 1 VSS VSS N18 L=1.8E-07 W=8E-07
M67 8 9 VSS VSS N18 L=1.8E-07 W=1.6E-06
M68 YX[1] 8 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M69 9 8 VSS VSS N18 L=1E-06 W=2.2E-07
M70 YCKX 8 YX[1] VSS N18 L=1.8E-07 W=1.25E-06
M71 29 5 23 VSS N18 L=1.8E-07 W=1E-06
M72 YX[1] 8 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M73 23 CLKX 9 VSS N18 L=1.8E-07 W=1.6E-06
M74 VSS 10 29 VSS N18 L=1.8E-07 W=1E-06
M75 YCKX 8 YX[1] VSS N18 L=1.8E-07 W=1.25E-06
M76 30 10 VSS VSS N18 L=1.8E-07 W=1E-06
M77 YX[3] 13 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M78 11 CLKX 24 VSS N18 L=1.8E-07 W=1.6E-06
M79 24 12 30 VSS N18 L=1.8E-07 W=1E-06
M80 YCKX 13 YX[3] VSS N18 L=1.8E-07 W=1.25E-06
M81 VSS 13 11 VSS N18 L=1E-06 W=2.2E-07
M82 YX[3] 13 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M83 VSS A[1] 5 VSS N18 L=1.8E-07 W=8E-07
M84 VSS 11 13 VSS N18 L=1.8E-07 W=1.6E-06
M85 YCKX 13 YX[3] VSS N18 L=1.8E-07 W=1.25E-06
M86 12 5 VSS VSS N18 L=1.8E-07 W=8E-07
M87 15 16 VSS VSS N18 L=1.8E-07 W=1.6E-06
M88 YX[2] 15 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M89 16 15 VSS VSS N18 L=1E-06 W=2.2E-07
M90 YCKX 15 YX[2] VSS N18 L=1.8E-07 W=1.25E-06
M91 31 12 27 VSS N18 L=1.8E-07 W=1E-06
M92 YX[2] 15 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M93 27 CLKX 16 VSS N18 L=1.8E-07 W=1.6E-06
M94 VSS 1 31 VSS N18 L=1.8E-07 W=1E-06
M95 YCKX 15 YX[2] VSS N18 L=1.8E-07 W=1.25E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_TP_CLKW_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_TP_CLKW_FLT CEN CLK DCTRCLK DCTRCLKX EMCLKB FB INTCLKX S[0] VDD VMINE VSS
M0 6 10 VDD VDD P18 L=1.8E-07 W=4E-06
M1 VDD 10 6 VDD P18 L=1.8E-07 W=4E-06
M2 3 6 VDD VDD P18 L=1.8E-07 W=2E-06
M3 VDD 6 3 VDD P18 L=1.8E-07 W=2E-06
M4 8 2 3 VDD P18 L=1.8E-07 W=2E-06
M5 3 2 8 VDD P18 L=1.8E-07 W=2E-06
M6 VDD S[0] 7 VDD P18 L=1.8E-07 W=8E-07
M7 1 7 VDD VDD P18 L=1.8E-07 W=1.2E-06
M8 2 1 VDD VDD P18 L=1.8E-07 W=1.2E-06
M9 8 1 29 VDD P18 L=1.8E-07 W=2E-06
M10 29 1 8 VDD P18 L=1.8E-07 W=2E-06
M11 29 6 VDD VDD P18 L=1.8E-07 W=2E-06
M12 VDD 5 29 VDD P18 L=1.8E-07 W=2E-06
M13 VDD 3 5 VDD P18 L=1.8E-07 W=2E-06
M14 EMCLKB 8 VDD VDD P18 L=1.8E-07 W=4E-06
M15 VDD 8 EMCLKB VDD P18 L=1.8E-07 W=4E-06
M16 11 FB VDD VDD P18 L=1.8E-07 W=1.2E-06
M17 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M18 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M19 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M20 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M21 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M22 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M23 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M24 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M25 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M26 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M27 VDD 15 9 VDD P18 L=1.8E-07 W=2.1E-06
M28 9 15 VDD VDD P18 L=1.8E-07 W=2.1E-06
M29 VDD 11 9 VDD P18 L=1.8E-07 W=2.1E-06
M30 9 11 VDD VDD P18 L=1.8E-07 W=2.1E-06
M31 VDD 15 35 VDD P18 L=1.8E-07 W=2E-06
M32 35 15 VDD VDD P18 L=1.8E-07 W=2E-06
M33 VDD 15 35 VDD P18 L=1.8E-07 W=2E-06
M34 35 15 VDD VDD P18 L=1.8E-07 W=2E-06
M35 VDD 15 35 VDD P18 L=1.8E-07 W=2E-06
M36 35 15 VDD VDD P18 L=1.8E-07 W=2E-06
M37 10 CLK 35 VDD P18 L=1.8E-07 W=2E-06
M38 35 CLK 10 VDD P18 L=1.8E-07 W=2E-06
M39 10 CLK 35 VDD P18 L=1.8E-07 W=2E-06
M40 35 CLK 10 VDD P18 L=1.8E-07 W=2E-06
M41 10 CLK 35 VDD P18 L=1.8E-07 W=2E-06
M42 35 CLK 10 VDD P18 L=1.8E-07 W=2E-06
M43 FB 6 VDD VDD P18 L=1.8E-07 W=2.4E-06
M44 VDD 6 FB VDD P18 L=1.8E-07 W=2.4E-06
M45 FB 6 VDD VDD P18 L=1.8E-07 W=2.4E-06
M46 17 10 VDD VDD P18 L=1.8E-07 W=9.95E-07
M47 VDD 10 17 VDD P18 L=1.8E-07 W=3.28E-06
M48 17 10 VDD VDD P18 L=1.8E-07 W=3.28E-06
M49 VDD 10 17 VDD P18 L=1.8E-07 W=3.28E-06
M50 17 10 VDD VDD P18 L=1.8E-07 W=3.28E-06
M51 15 VMINE VDD VDD P18 L=1.8E-07 W=2.8E-06
M52 42 CLK VDD VDD P18 L=1.8E-07 W=2E-06
M53 18 CEN 42 VDD P18 L=1.8E-07 W=2E-06
M54 43 16 VDD VDD P18 L=1.8E-07 W=2E-06
M55 19 CLK 43 VDD P18 L=1.8E-07 W=2E-06
M56 20 19 VDD VDD P18 L=1.8E-07 W=2E-06
M57 12 20 VDD VDD P18 L=1.8E-07 W=2E-06
M58 VDD 20 12 VDD P18 L=1.8E-07 W=2E-06
M59 12 20 VDD VDD P18 L=1.8E-07 W=2E-06
M60 VDD 16 18 VDD P18 L=1E-06 W=2.2E-07
M61 10 17 VDD VDD P18 L=1E-06 W=2.2E-07
M62 VDD CLK 21 VDD P18 L=1.8E-07 W=1.2E-06
M63 16 18 VDD VDD P18 L=1.8E-07 W=1.2E-06
M64 DCTRCLK 24 VDD VDD P18 L=1.8E-07 W=3.06E-06
M65 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=3.06E-06
M66 DCTRCLK 24 VDD VDD P18 L=1.8E-07 W=3.06E-06
M67 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=3.06E-06
M68 DCTRCLK 24 VDD VDD P18 L=1.8E-07 W=3.06E-06
M69 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=3.06E-06
M70 27 24 VDD VDD P18 L=1.8E-07 W=3E-06
M71 VDD 24 27 VDD P18 L=1.8E-07 W=3E-06
M72 24 17 38 VDD P18 L=1.8E-07 W=3.5E-06
M73 38 17 24 VDD P18 L=1.8E-07 W=3.5E-06
M74 VDD 26 38 VDD P18 L=1.8E-07 W=3.5E-06
M75 38 26 VDD VDD P18 L=1.8E-07 W=3.5E-06
M76 VDD 17 25 VDD P18 L=1.8E-07 W=5E-07
M77 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=1.66E-06
M78 VDD 17 INTCLKX VDD P18 L=1.8E-07 W=2.8E-06
M79 INTCLKX 17 VDD VDD P18 L=1.8E-07 W=2.8E-06
M80 VDD 17 INTCLKX VDD P18 L=1.8E-07 W=2.8E-06
M81 INTCLKX 17 VDD VDD P18 L=1.8E-07 W=2.8E-06
M82 VDD 17 INTCLKX VDD P18 L=1.8E-07 W=2.8E-06
M83 VDD 25 26 VDD P18 L=1.8E-07 W=5E-07
M84 DCTRCLKX 27 VDD VDD P18 L=1.8E-07 W=6.67E-06
M85 VDD 27 DCTRCLKX VDD P18 L=1.8E-07 W=6.67E-06
M86 DCTRCLKX 27 VDD VDD P18 L=1.8E-07 W=6.67E-06
M87 6 10 VSS VSS N18 L=1.8E-07 W=2E-06
M88 VSS 10 6 VSS N18 L=1.8E-07 W=2E-06
M89 3 6 VSS VSS N18 L=1.8E-07 W=2E-06
M90 VSS 6 3 VSS N18 L=1.8E-07 W=2E-06
M91 8 1 3 VSS N18 L=1.8E-07 W=2E-06
M92 3 1 8 VSS N18 L=1.8E-07 W=2E-06
M93 8 2 29 VSS N18 L=1.8E-07 W=2E-06
M94 29 2 8 VSS N18 L=1.8E-07 W=2E-06
M95 40 6 29 VSS N18 L=1.8E-07 W=2E-06
M96 VSS 5 40 VSS N18 L=1.8E-07 W=2E-06
M97 EMCLKB 8 VSS VSS N18 L=1.8E-07 W=2E-06
M98 VSS 8 EMCLKB VSS N18 L=1.8E-07 W=2E-06
M99 1 7 VSS VSS N18 L=1.8E-07 W=1.2E-06
M100 2 1 VSS VSS N18 L=1.8E-07 W=1.2E-06
M101 VSS 3 5 VSS N18 L=1.8E-07 W=1E-06
M102 VSS S[0] 7 VSS N18 L=1.8E-07 W=8E-07
M103 9 15 33 VSS N18 L=1.8E-07 W=2.1E-06
M104 33 15 9 VSS N18 L=1.8E-07 W=2.1E-06
M105 VSS 11 33 VSS N18 L=1.8E-07 W=2.1E-06
M106 33 11 VSS VSS N18 L=1.8E-07 W=2.1E-06
M107 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M108 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M109 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M110 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M111 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M112 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M113 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M114 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M115 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M116 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M117 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M118 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M119 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M120 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M121 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M122 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M123 11 FB VSS VSS N18 L=1.8E-07 W=1.2E-06
M124 VSS CLK 21 VSS N18 L=1.8E-07 W=1.2E-06
M125 41 21 VSS VSS N18 L=1.8E-07 W=2E-06
M126 18 CEN 41 VSS N18 L=1.8E-07 W=2E-06
M127 16 18 VSS VSS N18 L=1.8E-07 W=1.2E-06
M128 19 16 VSS VSS N18 L=1.8E-07 W=1E-06
M129 VSS CLK 19 VSS N18 L=1.8E-07 W=1E-06
M130 20 19 VSS VSS N18 L=1.8E-07 W=1E-06
M131 12 20 VSS VSS N18 L=1.8E-07 W=1.5E-06
M132 VSS 20 12 VSS N18 L=1.8E-07 W=1.5E-06
M133 VSS 10 17 VSS N18 L=1.8E-07 W=1.75E-06
M134 17 10 VSS VSS N18 L=1.8E-07 W=1.75E-06
M135 VSS 10 17 VSS N18 L=1.8E-07 W=1.75E-06
M136 17 10 VSS VSS N18 L=1.8E-07 W=1.75E-06
M137 10 17 VSS VSS N18 L=1E-06 W=2.2E-07
M138 18 16 VSS VSS N18 L=1E-06 W=2.2E-07
M139 15 VMINE VSS VSS N18 L=1.8E-07 W=1.4E-06
M140 24 17 VSS VSS N18 L=1.8E-07 W=3.5E-06
M141 VSS 17 24 VSS N18 L=1.8E-07 W=3.5E-06
M142 24 26 VSS VSS N18 L=1.8E-07 W=3.5E-06
M143 VSS 26 24 VSS N18 L=1.8E-07 W=3.5E-06
M144 VSS 24 DCTRCLK VSS N18 L=1.8E-07 W=3.335E-06
M145 DCTRCLK 24 VSS VSS N18 L=1.8E-07 W=3.335E-06
M146 VSS 24 DCTRCLK VSS N18 L=1.8E-07 W=3.335E-06
M147 27 24 VSS VSS N18 L=1.8E-07 W=3E-06
M148 VSS 24 27 VSS N18 L=1.8E-07 W=3E-06
M149 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=4.4E-06
M150 INTCLKX 17 VSS VSS N18 L=1.8E-07 W=4.4E-06
M151 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=4.4E-06
M152 INTCLKX 17 VSS VSS N18 L=1.8E-07 W=4.4E-06
M153 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=4.4E-06
M154 INTCLKX 17 VSS VSS N18 L=1.8E-07 W=3E-06
M155 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=3E-06
M156 VSS 25 26 VSS N18 L=1.8E-07 W=5E-07
M157 VSS 17 25 VSS N18 L=1.8E-07 W=5E-07
M158 DCTRCLKX 27 VSS VSS N18 L=1.8E-07 W=5E-06
M159 VSS 27 DCTRCLKX VSS N18 L=1.8E-07 W=5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_LOGIC_Y4_W_X64
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_LOGIC_Y4_W_X64 AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CENB CLKB
+DCTRCLK DCTRCLKX EMCLKB FB FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2]
+FCKXB[1] FCKXB[0] PXAB[3] PXAB[2] PXAB[1] PXAB[0] PXBB[1] PXBB[0] S[0] VDD
+VMINE VSS YXW[3] YXW[2] YXW[1] YXW[0]
XI0 AB[7] DCTRCLK DCTRCLKX PXBB[1] PXBB[0] VDD VSS RAM256_LEAFCELL_PX2_FLT
XPA AB[5] AB[6] DCTRCLK DCTRCLKX PXAB[3] PXAB[2] PXAB[1] PXAB[0] VDD VSS 
+ RAM256_LEAFCELL_PX4_FLT
XI37 AB[0] AB[1] DCTRCLK DCTRCLKX VDD VSS INTCLKXB YXW[3] YXW[2] YXW[1] YXW[0] 
+ RAM256_YPREDEC4_FLT
XFPRE AB[2] AB[3] AB[4] DCTRCLK DCTRCLKX FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] 
+ FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0] VDD VSS INTCLKXB RAM256_FPREDEC_FLT
XCLKDRV CENB CLKB DCTRCLK DCTRCLKX EMCLKB FB INTCLKXB S[0] VDD VMINE VSS 
+ RAM256_TP_CLKW_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_CLK_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_CLK_FLT ACTRCLK ACTRCLKX CEN CLK EMCLKA FB INTCLKX S[0] SACK1 SACK4
+VDD VMINE VSS
M0 4 VMINE VDD VDD P18 L=1.8E-07 W=2.8E-06
M1 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M2 7 2 VDD VDD P18 L=1.8E-07 W=4E-06
M3 ACTRCLKX ACTRCLK VDD VDD P18 L=1.8E-07 W=3.5E-06
M4 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M5 VDD 4 36 VDD P18 L=1.8E-07 W=2E-06
M6 VDD 2 7 VDD P18 L=1.8E-07 W=4E-06
M7 VDD ACTRCLK ACTRCLKX VDD P18 L=1.8E-07 W=3.5E-06
M8 VDD CLK 6 VDD P18 L=1.8E-07 W=1.2E-06
M9 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M10 36 4 VDD VDD P18 L=1.8E-07 W=2E-06
M11 ACTRCLKX ACTRCLK VDD VDD P18 L=1.8E-07 W=3.5E-06
M12 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M13 VDD 4 36 VDD P18 L=1.8E-07 W=2E-06
M14 47 CLK VDD VDD P18 L=1.8E-07 W=2E-06
M15 26 7 VDD VDD P18 L=1.8E-07 W=2E-06
M16 VDD ACTRCLK ACTRCLKX VDD P18 L=1.8E-07 W=3.5E-06
M17 10 CEN 47 VDD P18 L=1.8E-07 W=2E-06
M18 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M19 36 4 VDD VDD P18 L=1.8E-07 W=2E-06
M20 VDD 7 26 VDD P18 L=1.8E-07 W=2E-06
M21 ACTRCLK 11 VDD VDD P18 L=1.8E-07 W=3.5E-06
M22 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M23 VDD 4 36 VDD P18 L=1.8E-07 W=2E-06
M24 VDD 11 ACTRCLK VDD P18 L=1.8E-07 W=3.5E-06
M25 12 10 VDD VDD P18 L=1.8E-07 W=1.2E-06
M26 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M27 36 4 VDD VDD P18 L=1.8E-07 W=2E-06
M28 29 14 26 VDD P18 L=1.8E-07 W=2E-06
M29 ACTRCLK 11 VDD VDD P18 L=1.8E-07 W=3.5E-06
M30 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M31 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M32 2 CLK 36 VDD P18 L=1.8E-07 W=2E-06
M33 26 14 29 VDD P18 L=1.8E-07 W=2E-06
M34 VDD 11 ACTRCLK VDD P18 L=1.8E-07 W=3.5E-06
M35 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M36 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M37 36 CLK 2 VDD P18 L=1.8E-07 W=2E-06
M38 VDD 12 10 VDD P18 L=1E-06 W=2.2E-07
M39 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M40 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M41 2 CLK 36 VDD P18 L=1.8E-07 W=2E-06
M42 VDD S[0] 16 VDD P18 L=1.8E-07 W=8E-07
M43 11 9 38 VDD P18 L=1.8E-07 W=2.5E-06
M44 48 12 VDD VDD P18 L=1.8E-07 W=2E-06
M45 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M46 36 CLK 2 VDD P18 L=1.8E-07 W=2E-06
M47 38 9 11 VDD P18 L=1.8E-07 W=2.5E-06
M48 13 16 VDD VDD P18 L=1.8E-07 W=1.2E-06
M49 19 CLK 48 VDD P18 L=1.8E-07 W=2E-06
M50 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M51 2 CLK 36 VDD P18 L=1.8E-07 W=2E-06
M52 VDD 18 38 VDD P18 L=1.8E-07 W=2.5E-06
M53 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M54 36 CLK 2 VDD P18 L=1.8E-07 W=2E-06
M55 38 18 VDD VDD P18 L=1.8E-07 W=2.5E-06
M56 14 13 VDD VDD P18 L=1.8E-07 W=1.2E-06
M57 21 19 VDD VDD P18 L=1.8E-07 W=2E-06
M58 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M59 SACK1 9 VDD VDD P18 L=1.8E-07 W=1.86E-06
M60 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M61 29 13 39 VDD P18 L=1.8E-07 W=2E-06
M62 FB 7 VDD VDD P18 L=1.8E-07 W=2.4E-06
M63 VDD 9 SACK1 VDD P18 L=1.8E-07 W=3.035E-06
M64 20 21 VDD VDD P18 L=1.8E-07 W=2E-06
M65 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M66 VDD 22 18 VDD P18 L=1.8E-07 W=5E-07
M67 VDD 9 22 VDD P18 L=1.8E-07 W=5E-07
M68 39 13 29 VDD P18 L=1.8E-07 W=2E-06
M69 VDD 7 FB VDD P18 L=1.8E-07 W=2.4E-06
M70 SACK1 9 VDD VDD P18 L=1.8E-07 W=3.035E-06
M71 VDD 21 20 VDD P18 L=1.8E-07 W=2E-06
M72 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M73 FB 7 VDD VDD P18 L=1.8E-07 W=2.4E-06
M74 VDD 9 SACK1 VDD P18 L=1.8E-07 W=3.035E-06
M75 20 21 VDD VDD P18 L=1.8E-07 W=2E-06
M76 39 7 VDD VDD P18 L=1.8E-07 W=2E-06
M77 SACK1 9 VDD VDD P18 L=1.8E-07 W=3.035E-06
M78 24 9 VDD VDD P18 L=1.8E-07 W=5E-07
M79 28 24 VDD VDD P18 L=1.8E-07 W=5E-07
M80 30 FB VDD VDD P18 L=1.8E-07 W=1.2E-06
M81 2 9 VDD VDD P18 L=1E-06 W=2.2E-07
M82 VDD 25 39 VDD P18 L=1.8E-07 W=2E-06
M83 9 2 VDD VDD P18 L=1.8E-07 W=9.95E-07
M84 VDD 27 SACK4 VDD P18 L=1.8E-07 W=2.8E-06
M85 VDD 26 25 VDD P18 L=1.8E-07 W=2E-06
M86 VDD 4 17 VDD P18 L=1.8E-07 W=2.1E-06
M87 VDD 2 9 VDD P18 L=1.8E-07 W=3.28E-06
M88 43 9 27 VDD P18 L=1.8E-07 W=3E-06
M89 SACK4 27 VDD VDD P18 L=1.8E-07 W=2.8E-06
M90 17 4 VDD VDD P18 L=1.8E-07 W=2.1E-06
M91 9 2 VDD VDD P18 L=1.8E-07 W=3.28E-06
M92 VDD 28 43 VDD P18 L=1.8E-07 W=3E-06
M93 VDD 27 SACK4 VDD P18 L=1.8E-07 W=2.8E-06
M94 EMCLKA 29 VDD VDD P18 L=1.8E-07 W=4E-06
M95 VDD 30 17 VDD P18 L=1.8E-07 W=2.1E-06
M96 VDD 2 9 VDD P18 L=1.8E-07 W=3.28E-06
M97 43 28 VDD VDD P18 L=1.8E-07 W=3E-06
M98 SACK4 27 VDD VDD P18 L=1.8E-07 W=2.8E-06
M99 VDD 29 EMCLKA VDD P18 L=1.8E-07 W=4E-06
M100 17 30 VDD VDD P18 L=1.8E-07 W=2.1E-06
M101 9 2 VDD VDD P18 L=1.8E-07 W=3.28E-06
M102 27 9 43 VDD P18 L=1.8E-07 W=3E-06
M103 VDD 27 SACK4 VDD P18 L=1.8E-07 W=2.8E-06
M104 4 VMINE VSS VSS N18 L=1.8E-07 W=1.4E-06
M105 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M106 7 2 VSS VSS N18 L=1.8E-07 W=2E-06
M107 ACTRCLKX ACTRCLK VSS VSS N18 L=1.8E-07 W=1.75E-06
M108 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M109 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M110 VSS 2 7 VSS N18 L=1.8E-07 W=2E-06
M111 VSS ACTRCLK ACTRCLKX VSS N18 L=1.8E-07 W=1.75E-06
M112 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M113 VSS CLK 6 VSS N18 L=1.8E-07 W=1.2E-06
M114 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M115 ACTRCLKX ACTRCLK VSS VSS N18 L=1.8E-07 W=1.75E-06
M116 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M117 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M118 45 6 VSS VSS N18 L=1.8E-07 W=2E-06
M119 26 7 VSS VSS N18 L=1.8E-07 W=2E-06
M120 VSS ACTRCLK ACTRCLKX VSS N18 L=1.8E-07 W=1.75E-06
M121 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M122 10 CEN 45 VSS N18 L=1.8E-07 W=2E-06
M123 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M124 VSS 7 26 VSS N18 L=1.8E-07 W=2E-06
M125 ACTRCLK 11 VSS VSS N18 L=1.8E-07 W=1.75E-06
M126 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M127 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M128 VSS 11 ACTRCLK VSS N18 L=1.8E-07 W=1.75E-06
M129 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M130 12 10 VSS VSS N18 L=1.8E-07 W=1.2E-06
M131 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M132 29 13 26 VSS N18 L=1.8E-07 W=2E-06
M133 ACTRCLK 11 VSS VSS N18 L=1.8E-07 W=1.75E-06
M134 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M135 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M136 26 13 29 VSS N18 L=1.8E-07 W=2E-06
M137 VSS 11 ACTRCLK VSS N18 L=1.8E-07 W=1.75E-06
M138 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M139 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M140 10 12 VSS VSS N18 L=1E-06 W=2.2E-07
M141 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M142 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M143 VSS S[0] 16 VSS N18 L=1.8E-07 W=8E-07
M144 11 9 VSS VSS N18 L=1.8E-07 W=2.5E-06
M145 19 12 VSS VSS N18 L=1.8E-07 W=1E-06
M146 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M147 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M148 VSS 9 11 VSS N18 L=1.8E-07 W=2.5E-06
M149 13 16 VSS VSS N18 L=1.8E-07 W=1.2E-06
M150 VSS CLK 19 VSS N18 L=1.8E-07 W=1E-06
M151 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M152 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M153 11 18 VSS VSS N18 L=1.8E-07 W=2.5E-06
M154 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M155 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=1.4E-06
M156 VSS 18 11 VSS N18 L=1.8E-07 W=2.5E-06
M157 14 13 VSS VSS N18 L=1.8E-07 W=1.2E-06
M158 21 19 VSS VSS N18 L=1.8E-07 W=1E-06
M159 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M160 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=1.4E-06
M161 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M162 29 14 39 VSS N18 L=1.8E-07 W=2E-06
M163 20 21 VSS VSS N18 L=1.8E-07 W=1.5E-06
M164 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M165 VSS 22 18 VSS N18 L=1.8E-07 W=5E-07
M166 VSS 9 22 VSS N18 L=1.8E-07 W=5E-07
M167 39 14 29 VSS N18 L=1.8E-07 W=2E-06
M168 SACK1 9 VSS VSS N18 L=1.8E-07 W=1.75E-06
M169 VSS 21 20 VSS N18 L=1.8E-07 W=1.5E-06
M170 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M171 VSS 9 SACK1 VSS N18 L=1.8E-07 W=1.75E-06
M172 2 9 VSS VSS N18 L=1E-06 W=2.2E-07
M173 46 7 39 VSS N18 L=1.8E-07 W=2E-06
M174 SACK1 9 VSS VSS N18 L=1.8E-07 W=1.75E-06
M175 24 9 VSS VSS N18 L=1.8E-07 W=5E-07
M176 28 24 VSS VSS N18 L=1.8E-07 W=5E-07
M177 30 FB VSS VSS N18 L=1.8E-07 W=1.2E-06
M178 VSS 25 46 VSS N18 L=1.8E-07 W=2E-06
M179 VSS 9 SACK1 VSS N18 L=1.8E-07 W=1.75E-06
M180 VSS 26 25 VSS N18 L=1.8E-07 W=1E-06
M181 17 4 42 VSS N18 L=1.8E-07 W=2.1E-06
M182 VSS 2 9 VSS N18 L=1.8E-07 W=1.75E-06
M183 27 9 VSS VSS N18 L=1.8E-07 W=1.5E-06
M184 SACK4 27 VSS VSS N18 L=1.8E-07 W=1.75E-06
M185 42 4 17 VSS N18 L=1.8E-07 W=2.1E-06
M186 9 2 VSS VSS N18 L=1.8E-07 W=1.75E-06
M187 VSS 28 27 VSS N18 L=1.8E-07 W=1.5E-06
M188 VSS 27 SACK4 VSS N18 L=1.8E-07 W=1.75E-06
M189 EMCLKA 29 VSS VSS N18 L=1.8E-07 W=2E-06
M190 VSS 30 42 VSS N18 L=1.8E-07 W=2.1E-06
M191 VSS 2 9 VSS N18 L=1.8E-07 W=1.75E-06
M192 27 28 VSS VSS N18 L=1.8E-07 W=1.5E-06
M193 SACK4 27 VSS VSS N18 L=1.8E-07 W=1.75E-06
M194 VSS 29 EMCLKA VSS N18 L=1.8E-07 W=2E-06
M195 42 30 VSS VSS N18 L=1.8E-07 W=2.1E-06
M196 9 2 VSS VSS N18 L=1.8E-07 W=1.75E-06
M197 VSS 9 27 VSS N18 L=1.8E-07 W=1.5E-06
M198 VSS 27 SACK4 VSS N18 L=1.8E-07 W=1.75E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_LOGIC_Y4_R_X64
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_LOGIC_Y4_R_X64 AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] CENA CLKA
+EMCLKA FB FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0]
+PXAA[3] PXAA[2] PXAA[1] PXAA[0] PXBA[1] PXBA[0] S[0] SACK1 SACK4 VDD
+VMINE VSS YXR[3] YXR[2] YXR[1] YXR[0]
XI3 AA[7] ACTRCLK ACTRCLKX PXBA[1] PXBA[0] VDD VSS RAM256_LEAFCELL_PX2_FLT
XFPRE AA[2] AA[3] AA[4] ACTRCLK ACTRCLKX FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] 
+ FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0] VDD VSS INTCLKXA RAM256_FPREDEC_FLT
XPXA4A AA[5] AA[6] ACTRCLK ACTRCLKX PXAA[3] PXAA[2] PXAA[1] PXAA[0] VDD VSS 
+ RAM256_LEAFCELL_PX4_FLT
XI2 AA[0] AA[1] ACTRCLK ACTRCLKX VDD VSS INTCLKXA YXR[3] YXR[2] YXR[1] YXR[0] 
+ RAM256_YPREDEC4_FLT
XCLKDRV ACTRCLK ACTRCLKX CENA CLKA EMCLKA FB INTCLKXA S[0] SACK1 SACK4 VDD 
+ VMINE VSS RAM256_CLK_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_XDEC_FLT
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_XDEC_FLT FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA PXB
+PXC VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
M0 6 4 VDD VDD P18 L=1.8E-07 W=1E-06
M1 VDD 4 6 VDD P18 L=1.8E-07 W=1E-06
M2 4 5 VDD VDD P18 L=1.8E-07 W=1.5E-06
M3 VDD 5 4 VDD P18 L=1.8E-07 W=1.5E-06
M4 VDD PXA 5 VDD P18 L=1.8E-07 W=1E-06
M5 5 PXB VDD VDD P18 L=1.8E-07 W=1E-06
M6 VDD PXC 5 VDD P18 L=1.8E-07 W=1E-06
M7 VDD 4 7 VDD P18 L=1.8E-07 W=1E-06
M8 8 4 VDD VDD P18 L=1.8E-07 W=1E-06
M9 VDD 4 9 VDD P18 L=1.8E-07 W=1E-06
M10 10 4 VDD VDD P18 L=1.8E-07 W=1E-06
M11 VDD 4 11 VDD P18 L=1.8E-07 W=1E-06
M12 12 4 VDD VDD P18 L=1.8E-07 W=1E-06
M13 VDD 4 13 VDD P18 L=1.8E-07 W=1E-06
M14 14 4 VDD VDD P18 L=1.8E-07 W=1E-06
M15 7 6 FCKX[0] VDD P18 L=1.8E-07 W=8E-07
M16 FCKX[1] 6 8 VDD P18 L=1.8E-07 W=8E-07
M17 9 6 FCKX[2] VDD P18 L=1.8E-07 W=8E-07
M18 FCKX[3] 6 10 VDD P18 L=1.8E-07 W=8E-07
M19 11 6 FCKX[4] VDD P18 L=1.8E-07 W=8E-07
M20 FCKX[5] 6 12 VDD P18 L=1.8E-07 W=8E-07
M21 13 6 FCKX[6] VDD P18 L=1.8E-07 W=8E-07
M22 FCKX[7] 6 14 VDD P18 L=1.8E-07 W=8E-07
M23 15 7 VDD VDD P18 L=1.8E-07 W=8E-07
M24 VDD 7 15 VDD P18 L=1.8E-07 W=8E-07
M25 16 8 VDD VDD P18 L=1.8E-07 W=8E-07
M26 VDD 8 16 VDD P18 L=1.8E-07 W=8E-07
M27 17 9 VDD VDD P18 L=1.8E-07 W=8E-07
M28 VDD 9 17 VDD P18 L=1.8E-07 W=8E-07
M29 18 10 VDD VDD P18 L=1.8E-07 W=8E-07
M30 VDD 10 18 VDD P18 L=1.8E-07 W=8E-07
M31 19 11 VDD VDD P18 L=1.8E-07 W=8E-07
M32 VDD 11 19 VDD P18 L=1.8E-07 W=8E-07
M33 20 12 VDD VDD P18 L=1.8E-07 W=8E-07
M34 VDD 12 20 VDD P18 L=1.8E-07 W=8E-07
M35 21 13 VDD VDD P18 L=1.8E-07 W=8E-07
M36 VDD 13 21 VDD P18 L=1.8E-07 W=8E-07
M37 22 14 VDD VDD P18 L=1.8E-07 W=8E-07
M38 VDD 14 22 VDD P18 L=1.8E-07 W=8E-07
M39 23 15 VDD VDD P18 L=1.8E-07 W=2E-06
M40 VDD 15 23 VDD P18 L=1.8E-07 W=2E-06
M41 24 16 VDD VDD P18 L=1.8E-07 W=2E-06
M42 VDD 16 24 VDD P18 L=1.8E-07 W=2E-06
M43 25 17 VDD VDD P18 L=1.8E-07 W=2E-06
M44 VDD 17 25 VDD P18 L=1.8E-07 W=2E-06
M45 26 18 VDD VDD P18 L=1.8E-07 W=2E-06
M46 VDD 18 26 VDD P18 L=1.8E-07 W=2E-06
M47 27 19 VDD VDD P18 L=1.8E-07 W=2E-06
M48 VDD 19 27 VDD P18 L=1.8E-07 W=2E-06
M49 28 20 VDD VDD P18 L=1.8E-07 W=2E-06
M50 VDD 20 28 VDD P18 L=1.8E-07 W=2E-06
M51 29 21 VDD VDD P18 L=1.8E-07 W=2E-06
M52 VDD 21 29 VDD P18 L=1.8E-07 W=2E-06
M53 30 22 VDD VDD P18 L=1.8E-07 W=2E-06
M54 VDD 22 30 VDD P18 L=1.8E-07 W=2E-06
M55 WL[0] 23 VDD VDD P18 L=1.8E-07 W=7E-06
M56 VDD 23 WL[0] VDD P18 L=1.8E-07 W=7E-06
M57 WL[1] 24 VDD VDD P18 L=1.8E-07 W=7E-06
M58 VDD 24 WL[1] VDD P18 L=1.8E-07 W=7E-06
M59 WL[2] 25 VDD VDD P18 L=1.8E-07 W=7E-06
M60 VDD 25 WL[2] VDD P18 L=1.8E-07 W=7E-06
M61 WL[3] 26 VDD VDD P18 L=1.8E-07 W=7E-06
M62 VDD 26 WL[3] VDD P18 L=1.8E-07 W=7E-06
M63 WL[4] 27 VDD VDD P18 L=1.8E-07 W=7E-06
M64 VDD 27 WL[4] VDD P18 L=1.8E-07 W=7E-06
M65 WL[5] 28 VDD VDD P18 L=1.8E-07 W=7E-06
M66 VDD 28 WL[5] VDD P18 L=1.8E-07 W=7E-06
M67 WL[6] 29 VDD VDD P18 L=1.8E-07 W=7E-06
M68 VDD 29 WL[6] VDD P18 L=1.8E-07 W=7E-06
M69 WL[7] 30 VDD VDD P18 L=1.8E-07 W=7E-06
M70 VDD 30 WL[7] VDD P18 L=1.8E-07 W=7E-06
M71 78 PXA 5 VSS N18 L=1.8E-07 W=1.6E-06
M72 79 PXB 78 VSS N18 L=1.8E-07 W=1.6E-06
M73 VSS PXC 79 VSS N18 L=1.8E-07 W=1.6E-06
M74 6 4 VSS VSS N18 L=1.8E-07 W=1E-06
M75 VSS 4 6 VSS N18 L=1.8E-07 W=1E-06
M76 4 5 VSS VSS N18 L=1.8E-07 W=1E-06
M77 VSS 5 4 VSS N18 L=1.8E-07 W=1E-06
M78 7 4 FCKX[0] VSS N18 L=1.8E-07 W=1E-06
M79 FCKX[1] 4 8 VSS N18 L=1.8E-07 W=1E-06
M80 9 4 FCKX[2] VSS N18 L=1.8E-07 W=1E-06
M81 FCKX[3] 4 10 VSS N18 L=1.8E-07 W=1E-06
M82 11 4 FCKX[4] VSS N18 L=1.8E-07 W=1E-06
M83 FCKX[5] 4 12 VSS N18 L=1.8E-07 W=1E-06
M84 13 4 FCKX[6] VSS N18 L=1.8E-07 W=1E-06
M85 FCKX[7] 4 14 VSS N18 L=1.8E-07 W=1E-06
M86 15 7 VSS VSS N18 L=1.8E-07 W=4E-07
M87 VSS 7 15 VSS N18 L=1.8E-07 W=4E-07
M88 16 8 VSS VSS N18 L=1.8E-07 W=4E-07
M89 VSS 8 16 VSS N18 L=1.8E-07 W=4E-07
M90 17 9 VSS VSS N18 L=1.8E-07 W=4E-07
M91 VSS 9 17 VSS N18 L=1.8E-07 W=4E-07
M92 18 10 VSS VSS N18 L=1.8E-07 W=4E-07
M93 VSS 10 18 VSS N18 L=1.8E-07 W=4E-07
M94 19 11 VSS VSS N18 L=1.8E-07 W=4E-07
M95 VSS 11 19 VSS N18 L=1.8E-07 W=4E-07
M96 20 12 VSS VSS N18 L=1.8E-07 W=4E-07
M97 VSS 12 20 VSS N18 L=1.8E-07 W=4E-07
M98 21 13 VSS VSS N18 L=1.8E-07 W=4E-07
M99 VSS 13 21 VSS N18 L=1.8E-07 W=4E-07
M100 22 14 VSS VSS N18 L=1.8E-07 W=4E-07
M101 VSS 14 22 VSS N18 L=1.8E-07 W=4E-07
M102 23 15 VSS VSS N18 L=1.8E-07 W=1.2E-06
M103 VSS 15 23 VSS N18 L=1.8E-07 W=1.2E-06
M104 24 16 VSS VSS N18 L=1.8E-07 W=1.2E-06
M105 VSS 16 24 VSS N18 L=1.8E-07 W=1.2E-06
M106 25 17 VSS VSS N18 L=1.8E-07 W=1.2E-06
M107 VSS 17 25 VSS N18 L=1.8E-07 W=1.2E-06
M108 26 18 VSS VSS N18 L=1.8E-07 W=1.2E-06
M109 VSS 18 26 VSS N18 L=1.8E-07 W=1.2E-06
M110 27 19 VSS VSS N18 L=1.8E-07 W=1.2E-06
M111 VSS 19 27 VSS N18 L=1.8E-07 W=1.2E-06
M112 28 20 VSS VSS N18 L=1.8E-07 W=1.2E-06
M113 VSS 20 28 VSS N18 L=1.8E-07 W=1.2E-06
M114 29 21 VSS VSS N18 L=1.8E-07 W=1.2E-06
M115 VSS 21 29 VSS N18 L=1.8E-07 W=1.2E-06
M116 30 22 VSS VSS N18 L=1.8E-07 W=1.2E-06
M117 VSS 22 30 VSS N18 L=1.8E-07 W=1.2E-06
M118 WL[0] 23 VSS VSS N18 L=1.8E-07 W=3.5E-06
M119 VSS 23 WL[0] VSS N18 L=1.8E-07 W=3.5E-06
M120 WL[1] 24 VSS VSS N18 L=1.8E-07 W=3.5E-06
M121 VSS 24 WL[1] VSS N18 L=1.8E-07 W=3.5E-06
M122 WL[2] 25 VSS VSS N18 L=1.8E-07 W=3.5E-06
M123 VSS 25 WL[2] VSS N18 L=1.8E-07 W=3.5E-06
M124 WL[3] 26 VSS VSS N18 L=1.8E-07 W=3.5E-06
M125 VSS 26 WL[3] VSS N18 L=1.8E-07 W=3.5E-06
M126 WL[4] 27 VSS VSS N18 L=1.8E-07 W=3.5E-06
M127 VSS 27 WL[4] VSS N18 L=1.8E-07 W=3.5E-06
M128 WL[5] 28 VSS VSS N18 L=1.8E-07 W=3.5E-06
M129 VSS 28 WL[5] VSS N18 L=1.8E-07 W=3.5E-06
M130 WL[6] 29 VSS VSS N18 L=1.8E-07 W=3.5E-06
M131 VSS 29 WL[6] VSS N18 L=1.8E-07 W=3.5E-06
M132 WL[7] 30 VSS VSS N18 L=1.8E-07 W=3.5E-06
M133 VSS 30 WL[7] VSS N18 L=1.8E-07 W=3.5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256_XDEC8
* View Name:    schematic
************************************************************************

.SUBCKT RAM256_XDEC8 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2]
+PXA[1] PXA[0] PXB[1] PXB[0] PXC[0] VDD VSS WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
XI0 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[0] VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] RAM256_XDEC_FLT
XI1 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[0] VDD VSS WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] RAM256_XDEC_FLT
XI2 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[0] VDD VSS WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] RAM256_XDEC_FLT
XI3 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[0] VDD VSS WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] RAM256_XDEC_FLT
XI4 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[0] VDD VSS WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] RAM256_XDEC_FLT
XI5 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[0] VDD VSS WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] RAM256_XDEC_FLT
XI6 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[0] VDD VSS WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] RAM256_XDEC_FLT
XI7 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[0] VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0] RAM256_XDEC_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    RAM256
* View Name:    schematic
************************************************************************

.SUBCKT RAM256 AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] AB[7] AB[6]
+AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CENA CENB CLKA CLKB
+DB[23] DB[22] DB[21] DB[20] DB[19] DB[18] DB[17] DB[16] DB[15] DB[14]
+DB[13] DB[12] DB[11] DB[10] DB[9] DB[8] DB[7] DB[6] DB[5] DB[4]
+DB[3] DB[2] DB[1] DB[0] QA[23] QA[22] QA[21] QA[20] QA[19] QA[18]
+QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] QA[11] QA[10] QA[9] QA[8]
+QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] VDD VSS
XI0 DCTRCLK DCTRCLKX DB[23] DB[22] DB[21] DB[20] DB[19] DB[18] DB[17] DB[16]
+DB[15] DB[14] DB[13] DB[12] DBLA QA[23] QA[22] QA[21] QA[20] QA[19]
+QA[18] QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] SACK1 SACK4 STWLA
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXR[3] YXR[2] YXR[1] YXR[0] YXW[3] YXW[2] YXW[1] YXW[0] RAM256_ARRAY_X64Y4D12_RIGHT
XI1 DCTRCLK DCTRCLKX DB[11] DB[10] DB[9] DB[8] DB[7] DB[6] DB[5] DB[4]
+DB[3] DB[2] DB[1] DB[0] DBLB QA[11] QA[10] QA[9] QA[8] QA[7]
+QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] SACK1 SACK4 STWLA
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+YXR[3] YXR[2] YXR[1] YXR[0] YXW[3] YXW[2] YXW[1] YXW[0] RAM256_ARRAY_X64Y4D12_LEFT
XI2 DBLA EMCLKA VSS VDD STWLA VDD VSS RAM256_SOP_FLT
XI3 DBLB EMCLKB VSS VDD VDD VSS RAM256_SOP_W_FLT
XI4 AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CENB CLKB
+DCTRCLK DCTRCLKX EMCLKB DBLB FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2]
+FCKXB[1] FCKXB[0] PXAB[3] PXAB[2] PXAB[1] PXAB[0] PXBB[1] PXBB[0] VSS VDD
+VSS VSS YXW[3] YXW[2] YXW[1] YXW[0] RAM256_LOGIC_Y4_W_X64
XI5 AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] CENA CLKA
+EMCLKA DBLA FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0]
+PXAA[3] PXAA[2] PXAA[1] PXAA[0] PXBA[1] PXBA[0] VSS SACK1 SACK4 VDD
+VSS VSS YXR[3] YXR[2] YXR[1] YXR[0] RAM256_LOGIC_Y4_R_X64
XI6 FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0] PXAB[3] PXAB[2]
+PXAB[1] PXAB[0] PXBB[1] PXBB[0] VDD VDD VSS WLB[63] WLB[62] WLB[61]
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51]
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41]
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31]
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21]
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11]
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1]
+WLB[0] RAM256_XDEC8
XI7 FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0] PXAA[3] PXAA[2]
+PXAA[1] PXAA[0] PXBA[1] PXBA[0] VDD VDD VSS WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41]
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31]
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1]
+WLA[0] RAM256_XDEC8
.ENDS
