#     Copyright (c) 2022 SMIC                                                       
#     Filename:      RAM128.lef                                                   
#     IP code:       S018RF2P                                                         
#     Version:       0.2.b                                                        
#     CreateDate:    Mon Oct 31 21:44:19 CST 2022                                                     
                    
#    LEF for 2-PORT Register File                                                               
#    SMIC 0.18um G Logic Process                                                       
#    Configuration: -instname RAM128 -rows 32 -bits 24 -mux 4  



# DISCLAIMER                                                                           #
#                                                                                      #  
#   SMIC hereby provides the quality information to you but makes no claims,           #
# promises or guarantees about the accuracy, completeness, or adequacy of the          #
# information herein. The information contained herein is provided on an "AS IS"       #
# basis without any warranty, and SMIC assumes no obligation to provide support        #
# of any kind or otherwise maintain the information.                                   #  
#   SMIC disclaims any representation that the information does not infringe any       #
# intellectual property rights or proprietary rights of any third parties. SMIC        #
# makes no other warranty, whether express, implied or statutory as to any             #
# matter whatsoever, including but not limited to the accuracy or sufficiency of       #
# any information or the merchantability and fitness for a particular purpose.         #
# Neither SMIC nor any of its representatives shall be liable for any cause of         #
# action incurred to connect to this service.                                          #  
#                                                                                      #
# STATEMENT OF USE AND CONFIDENTIALITY                                                 #  
#                                                                                      #  
#   The following/attached material contains confidential and proprietary              #  
# information of SMIC. This material is based upon information which SMIC              #  
# considers reliable, but SMIC neither represents nor warrants that such               #
# information is accurate or complete, and it must not be relied upon as such.         #
# This information was prepared for informational purposes and is for the use          #
# by SMIC's customer only. SMIC reserves the right to make changes in the              #  
# information at any time without notice.                                              #  
#   No part of this information may be reproduced, transmitted, transcribed,           #  
# stored in a retrieval system, or translated into any human or computer               # 
# language, in any form or by any means, electronic, mechanical, magnetic,             #  
# optical, chemical, manual, or otherwise, without the prior written consent of        #
# SMIC. Any unauthorized use or disclosure of this material is strictly                #  
# prohibited and may be unlawful. By accepting this material, the receiving            #  
# party shall be deemed to have acknowledged, accepted, and agreed to be bound         #
# by the foregoing limitations and restrictions. Thank you.                            #  
#                                                                                      #  


MACRO RAM128
CLASS BLOCK ;
ORIGIN 0 0 ;
SIZE 665.14 BY 103.4 ;
SYMMETRY X Y R90 ;

PIN QA[11]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 8.905 102.76 9.975 103.4 ;
LAYER METAL2 ;
RECT 8.905 102.76 9.975 103.4 ;
LAYER METAL3 ;
RECT 8.905 102.76 9.975 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[11]

PIN DB[11]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL2 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL3 ;
RECT 18.725 0.0 19.795 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[11]

PIN QA[10]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 32.145 102.76 33.215 103.4 ;
LAYER METAL2 ;
RECT 32.145 102.76 33.215 103.4 ;
LAYER METAL3 ;
RECT 32.145 102.76 33.215 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[10]

PIN DB[10]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL2 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL3 ;
RECT 41.965 0.0 43.035 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[10]

PIN QA[9]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 55.385 102.76 56.455 103.4 ;
LAYER METAL2 ;
RECT 55.385 102.76 56.455 103.4 ;
LAYER METAL3 ;
RECT 55.385 102.76 56.455 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[9]

PIN DB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL2 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL3 ;
RECT 65.205 0.0 66.275 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[9]

PIN QA[8]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 78.625 102.76 79.695 103.4 ;
LAYER METAL2 ;
RECT 78.625 102.76 79.695 103.4 ;
LAYER METAL3 ;
RECT 78.625 102.76 79.695 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[8]

PIN DB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL2 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL3 ;
RECT 88.445 0.0 89.515 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[8]

PIN QA[7]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 101.865 102.76 102.935 103.4 ;
LAYER METAL2 ;
RECT 101.865 102.76 102.935 103.4 ;
LAYER METAL3 ;
RECT 101.865 102.76 102.935 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[7]

PIN DB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL2 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL3 ;
RECT 111.685 0.0 112.755 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[7]

PIN QA[6]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 125.105 102.76 126.175 103.4 ;
LAYER METAL2 ;
RECT 125.105 102.76 126.175 103.4 ;
LAYER METAL3 ;
RECT 125.105 102.76 126.175 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[6]

PIN DB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL2 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL3 ;
RECT 134.925 0.0 135.995 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[6]

PIN QA[5]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 148.345 102.76 149.415 103.4 ;
LAYER METAL2 ;
RECT 148.345 102.76 149.415 103.4 ;
LAYER METAL3 ;
RECT 148.345 102.76 149.415 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[5]

PIN DB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL2 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL3 ;
RECT 158.165 0.0 159.235 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[5]

PIN QA[4]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 171.585 102.76 172.655 103.4 ;
LAYER METAL2 ;
RECT 171.585 102.76 172.655 103.4 ;
LAYER METAL3 ;
RECT 171.585 102.76 172.655 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[4]

PIN DB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL2 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL3 ;
RECT 181.405 0.0 182.475 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[4]

PIN QA[3]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 194.825 102.76 195.895 103.4 ;
LAYER METAL2 ;
RECT 194.825 102.76 195.895 103.4 ;
LAYER METAL3 ;
RECT 194.825 102.76 195.895 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[3]

PIN DB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL2 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL3 ;
RECT 204.645 0.0 205.715 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[3]

PIN QA[2]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 218.065 102.76 219.135 103.4 ;
LAYER METAL2 ;
RECT 218.065 102.76 219.135 103.4 ;
LAYER METAL3 ;
RECT 218.065 102.76 219.135 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[2]

PIN DB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL2 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL3 ;
RECT 227.885 0.0 228.955 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[2]

PIN QA[1]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 241.305 102.76 242.375 103.4 ;
LAYER METAL2 ;
RECT 241.305 102.76 242.375 103.4 ;
LAYER METAL3 ;
RECT 241.305 102.76 242.375 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[1]

PIN DB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL2 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL3 ;
RECT 251.125 0.0 252.195 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[1]

PIN QA[0]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 264.545 102.76 265.615 103.4 ;
LAYER METAL2 ;
RECT 264.545 102.76 265.615 103.4 ;
LAYER METAL3 ;
RECT 264.545 102.76 265.615 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[0]

PIN DB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL2 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL3 ;
RECT 274.365 0.0 275.435 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[0]

PIN CLKB
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL2 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL3 ;
RECT 297.105 0.0 297.605 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKB

PIN AA[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 297.655 102.76 298.905 103.4 ;
LAYER METAL2 ;
RECT 297.655 102.76 298.905 103.4 ;
LAYER METAL3 ;
RECT 297.655 102.76 298.905 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[0]

PIN AA[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 302.505 102.76 303.755 103.4 ;
LAYER METAL2 ;
RECT 302.505 102.76 303.755 103.4 ;
LAYER METAL3 ;
RECT 302.505 102.76 303.755 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[1]

PIN CENB
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL2 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL3 ;
RECT 306.72 0.0 307.22 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENB

PIN AA[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 312.875 102.76 314.525 103.4 ;
LAYER METAL2 ;
RECT 312.875 102.76 314.125 103.4 ;
LAYER METAL3 ;
RECT 312.875 102.76 314.125 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[4]

PIN AA[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 320.815 102.76 322.465 103.4 ;
LAYER METAL2 ;
RECT 320.815 102.76 322.065 103.4 ;
LAYER METAL3 ;
RECT 320.815 102.76 322.065 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[3]

PIN AB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 323.45 0.0 325.015 0.64 ;
LAYER METAL2 ;
RECT 323.765 0.0 325.015 0.64 ;
LAYER METAL3 ;
RECT 323.765 0.0 325.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[6]

PIN AA[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.755 102.76 330.405 103.4 ;
LAYER METAL2 ;
RECT 328.755 102.76 330.005 103.4 ;
LAYER METAL3 ;
RECT 328.755 102.76 330.005 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[2]

PIN AB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 329.21 0.0 330.775 0.64 ;
LAYER METAL2 ;
RECT 329.525 0.0 330.775 0.64 ;
LAYER METAL3 ;
RECT 329.525 0.0 330.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[5]

PIN AA[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.365 102.76 335.93 103.4 ;
LAYER METAL2 ;
RECT 334.365 102.76 335.615 103.4 ;
LAYER METAL3 ;
RECT 334.365 102.76 335.615 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[5]

PIN AB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.735 0.0 336.385 0.64 ;
LAYER METAL2 ;
RECT 335.135 0.0 336.385 0.64 ;
LAYER METAL3 ;
RECT 335.135 0.0 336.385 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[2]

PIN AA[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.125 102.76 341.69 103.4 ;
LAYER METAL2 ;
RECT 340.125 102.76 341.375 103.4 ;
LAYER METAL3 ;
RECT 340.125 102.76 341.375 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[6]

PIN AB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 342.675 0.0 344.325 0.64 ;
LAYER METAL2 ;
RECT 343.075 0.0 344.325 0.64 ;
LAYER METAL3 ;
RECT 343.075 0.0 344.325 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[3]

PIN AB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 350.615 0.0 352.265 0.64 ;
LAYER METAL2 ;
RECT 351.015 0.0 352.265 0.64 ;
LAYER METAL3 ;
RECT 351.015 0.0 352.265 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[4]

PIN CENA
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 359.765 102.33 360.265 103.4 ;
LAYER METAL2 ;
RECT 359.765 102.33 360.265 103.4 ;
LAYER METAL3 ;
RECT 359.765 102.33 360.265 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENA

PIN AB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 361.385 0.0 362.635 0.64 ;
LAYER METAL2 ;
RECT 361.385 0.0 362.635 0.64 ;
LAYER METAL3 ;
RECT 361.385 0.0 362.635 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[1]

PIN AB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 366.235 0.0 367.485 0.64 ;
LAYER METAL2 ;
RECT 366.235 0.0 367.485 0.64 ;
LAYER METAL3 ;
RECT 366.235 0.0 367.485 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[0]

PIN CLKA
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 369.17 102.33 369.67 103.4 ;
LAYER METAL2 ;
RECT 369.17 102.33 369.67 103.4 ;
LAYER METAL3 ;
RECT 369.17 102.33 369.67 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKA

PIN DB[12]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 389.705 0.0 390.775 0.64 ;
LAYER METAL2 ;
RECT 389.705 0.0 390.775 0.64 ;
LAYER METAL3 ;
RECT 389.705 0.0 390.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[12]

PIN QA[12]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 399.525 102.76 400.595 103.4 ;
LAYER METAL2 ;
RECT 399.525 102.76 400.595 103.4 ;
LAYER METAL3 ;
RECT 399.525 102.76 400.595 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[12]

PIN DB[13]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 412.945 0.0 414.015 0.64 ;
LAYER METAL2 ;
RECT 412.945 0.0 414.015 0.64 ;
LAYER METAL3 ;
RECT 412.945 0.0 414.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[13]

PIN QA[13]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 422.765 102.76 423.835 103.4 ;
LAYER METAL2 ;
RECT 422.765 102.76 423.835 103.4 ;
LAYER METAL3 ;
RECT 422.765 102.76 423.835 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[13]

PIN DB[14]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 436.185 0.0 437.255 0.64 ;
LAYER METAL2 ;
RECT 436.185 0.0 437.255 0.64 ;
LAYER METAL3 ;
RECT 436.185 0.0 437.255 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[14]

PIN QA[14]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 446.005 102.76 447.075 103.4 ;
LAYER METAL2 ;
RECT 446.005 102.76 447.075 103.4 ;
LAYER METAL3 ;
RECT 446.005 102.76 447.075 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[14]

PIN DB[15]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 459.425 0.0 460.495 0.64 ;
LAYER METAL2 ;
RECT 459.425 0.0 460.495 0.64 ;
LAYER METAL3 ;
RECT 459.425 0.0 460.495 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[15]

PIN QA[15]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 469.245 102.76 470.315 103.4 ;
LAYER METAL2 ;
RECT 469.245 102.76 470.315 103.4 ;
LAYER METAL3 ;
RECT 469.245 102.76 470.315 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[15]

PIN DB[16]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 482.665 0.0 483.735 0.64 ;
LAYER METAL2 ;
RECT 482.665 0.0 483.735 0.64 ;
LAYER METAL3 ;
RECT 482.665 0.0 483.735 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[16]

PIN QA[16]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 492.485 102.76 493.555 103.4 ;
LAYER METAL2 ;
RECT 492.485 102.76 493.555 103.4 ;
LAYER METAL3 ;
RECT 492.485 102.76 493.555 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[16]

PIN DB[17]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 505.905 0.0 506.975 0.64 ;
LAYER METAL2 ;
RECT 505.905 0.0 506.975 0.64 ;
LAYER METAL3 ;
RECT 505.905 0.0 506.975 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[17]

PIN QA[17]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 515.725 102.76 516.795 103.4 ;
LAYER METAL2 ;
RECT 515.725 102.76 516.795 103.4 ;
LAYER METAL3 ;
RECT 515.725 102.76 516.795 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[17]

PIN DB[18]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 529.145 0.0 530.215 0.64 ;
LAYER METAL2 ;
RECT 529.145 0.0 530.215 0.64 ;
LAYER METAL3 ;
RECT 529.145 0.0 530.215 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[18]

PIN QA[18]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 538.965 102.76 540.035 103.4 ;
LAYER METAL2 ;
RECT 538.965 102.76 540.035 103.4 ;
LAYER METAL3 ;
RECT 538.965 102.76 540.035 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[18]

PIN DB[19]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 552.385 0.0 553.455 0.64 ;
LAYER METAL2 ;
RECT 552.385 0.0 553.455 0.64 ;
LAYER METAL3 ;
RECT 552.385 0.0 553.455 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[19]

PIN QA[19]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 562.205 102.76 563.275 103.4 ;
LAYER METAL2 ;
RECT 562.205 102.76 563.275 103.4 ;
LAYER METAL3 ;
RECT 562.205 102.76 563.275 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[19]

PIN DB[20]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 575.625 0.0 576.695 0.64 ;
LAYER METAL2 ;
RECT 575.625 0.0 576.695 0.64 ;
LAYER METAL3 ;
RECT 575.625 0.0 576.695 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[20]

PIN QA[20]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 585.445 102.76 586.515 103.4 ;
LAYER METAL2 ;
RECT 585.445 102.76 586.515 103.4 ;
LAYER METAL3 ;
RECT 585.445 102.76 586.515 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[20]

PIN DB[21]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 598.865 0.0 599.935 0.64 ;
LAYER METAL2 ;
RECT 598.865 0.0 599.935 0.64 ;
LAYER METAL3 ;
RECT 598.865 0.0 599.935 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[21]

PIN QA[21]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 608.685 102.76 609.755 103.4 ;
LAYER METAL2 ;
RECT 608.685 102.76 609.755 103.4 ;
LAYER METAL3 ;
RECT 608.685 102.76 609.755 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[21]

PIN DB[22]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 622.105 0.0 623.175 0.64 ;
LAYER METAL2 ;
RECT 622.105 0.0 623.175 0.64 ;
LAYER METAL3 ;
RECT 622.105 0.0 623.175 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[22]

PIN QA[22]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 631.925 102.76 632.995 103.4 ;
LAYER METAL2 ;
RECT 631.925 102.76 632.995 103.4 ;
LAYER METAL3 ;
RECT 631.925 102.76 632.995 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[22]

PIN DB[23]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 645.345 0.0 646.415 0.64 ;
LAYER METAL2 ;
RECT 645.345 0.0 646.415 0.64 ;
LAYER METAL3 ;
RECT 645.345 0.0 646.415 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[23]

PIN QA[23]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 655.165 102.76 656.235 103.4 ;
LAYER METAL2 ;
RECT 655.165 102.76 656.235 103.4 ;
LAYER METAL3 ;
RECT 655.165 102.76 656.235 103.4 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[23]

PIN VSS
DIRECTION INOUT ;
USE GROUND ;
PORT
LAYER METAL4 ;
RECT 279.475 0.0 283.475 103.4 ;
LAYER METAL4 ;
RECT 290.475 0.0 294.475 103.4 ;
LAYER METAL4 ;
RECT 301.475 0.0 305.475 103.4 ;
LAYER METAL4 ;
RECT 312.475 0.0 316.475 103.4 ;
LAYER METAL4 ;
RECT 323.475 0.0 327.475 103.4 ;
LAYER METAL4 ;
RECT 337.665 0.0 341.665 103.4 ;
LAYER METAL4 ;
RECT 348.665 0.0 352.665 103.4 ;
LAYER METAL4 ;
RECT 359.665 0.0 363.665 103.4 ;
LAYER METAL4 ;
RECT 370.665 0.0 374.665 103.4 ;
LAYER METAL4 ;
RECT 381.665 0.0 385.665 103.4 ;
LAYER METAL4 ;
RECT 267.855 0.0 271.855 103.4 ;
LAYER METAL4 ;
RECT 256.235 0.0 260.235 103.4 ;
LAYER METAL4 ;
RECT 244.615 0.0 248.615 103.4 ;
LAYER METAL4 ;
RECT 232.995 0.0 236.995 103.4 ;
LAYER METAL4 ;
RECT 221.375 0.0 225.375 103.4 ;
LAYER METAL4 ;
RECT 209.755 0.0 213.755 103.4 ;
LAYER METAL4 ;
RECT 198.135 0.0 202.135 103.4 ;
LAYER METAL4 ;
RECT 186.515 0.0 190.515 103.4 ;
LAYER METAL4 ;
RECT 174.895 0.0 178.895 103.4 ;
LAYER METAL4 ;
RECT 163.275 0.0 167.275 103.4 ;
LAYER METAL4 ;
RECT 151.655 0.0 155.655 103.4 ;
LAYER METAL4 ;
RECT 140.035 0.0 144.035 103.4 ;
LAYER METAL4 ;
RECT 128.415 0.0 132.415 103.4 ;
LAYER METAL4 ;
RECT 116.795 0.0 120.795 103.4 ;
LAYER METAL4 ;
RECT 105.175 0.0 109.175 103.4 ;
LAYER METAL4 ;
RECT 93.555 0.0 97.555 103.4 ;
LAYER METAL4 ;
RECT 81.935 0.0 85.935 103.4 ;
LAYER METAL4 ;
RECT 70.315 0.0 74.315 103.4 ;
LAYER METAL4 ;
RECT 58.695 0.0 62.695 103.4 ;
LAYER METAL4 ;
RECT 47.075 0.0 51.075 103.4 ;
LAYER METAL4 ;
RECT 35.455 0.0 39.455 103.4 ;
LAYER METAL4 ;
RECT 23.835 0.0 27.835 103.4 ;
LAYER METAL4 ;
RECT 12.215 0.0 16.215 103.4 ;
LAYER METAL4 ;
RECT 0.595 0.0 4.595 103.4 ;
LAYER METAL4 ;
RECT 393.285 0.0 397.285 103.4 ;
LAYER METAL4 ;
RECT 404.905 0.0 408.905 103.4 ;
LAYER METAL4 ;
RECT 416.525 0.0 420.525 103.4 ;
LAYER METAL4 ;
RECT 428.145 0.0 432.145 103.4 ;
LAYER METAL4 ;
RECT 439.765 0.0 443.765 103.4 ;
LAYER METAL4 ;
RECT 451.385 0.0 455.385 103.4 ;
LAYER METAL4 ;
RECT 463.005 0.0 467.005 103.4 ;
LAYER METAL4 ;
RECT 474.625 0.0 478.625 103.4 ;
LAYER METAL4 ;
RECT 486.245 0.0 490.245 103.4 ;
LAYER METAL4 ;
RECT 497.865 0.0 501.865 103.4 ;
LAYER METAL4 ;
RECT 509.485 0.0 513.485 103.4 ;
LAYER METAL4 ;
RECT 521.105 0.0 525.105 103.4 ;
LAYER METAL4 ;
RECT 532.725 0.0 536.725 103.4 ;
LAYER METAL4 ;
RECT 544.345 0.0 548.345 103.4 ;
LAYER METAL4 ;
RECT 555.965 0.0 559.965 103.4 ;
LAYER METAL4 ;
RECT 567.585 0.0 571.585 103.4 ;
LAYER METAL4 ;
RECT 579.205 0.0 583.205 103.4 ;
LAYER METAL4 ;
RECT 590.825 0.0 594.825 103.4 ;
LAYER METAL4 ;
RECT 602.445 0.0 606.445 103.4 ;
LAYER METAL4 ;
RECT 614.065 0.0 618.065 103.4 ;
LAYER METAL4 ;
RECT 625.685 0.0 629.685 103.4 ;
LAYER METAL4 ;
RECT 637.305 0.0 641.305 103.4 ;
LAYER METAL4 ;
RECT 648.925 0.0 652.925 103.4 ;
LAYER METAL4 ;
RECT 660.545 0.0 664.545 103.4 ;
END
END VSS

PIN VDD
DIRECTION INOUT ;
USE POWER ;
PORT
LAYER METAL4 ;
RECT 284.975 0.0 288.975 103.4 ;
LAYER METAL4 ;
RECT 295.975 0.0 299.975 103.4 ;
LAYER METAL4 ;
RECT 306.975 0.0 310.975 103.4 ;
LAYER METAL4 ;
RECT 317.975 0.0 321.975 103.4 ;
LAYER METAL4 ;
RECT 343.165 0.0 347.165 103.4 ;
LAYER METAL4 ;
RECT 354.165 0.0 358.165 103.4 ;
LAYER METAL4 ;
RECT 365.165 0.0 369.165 103.4 ;
LAYER METAL4 ;
RECT 376.165 0.0 380.165 103.4 ;
LAYER METAL4 ;
RECT 273.665 0.0 277.665 103.4 ;
LAYER METAL4 ;
RECT 262.045 0.0 266.045 103.4 ;
LAYER METAL4 ;
RECT 250.425 0.0 254.425 103.4 ;
LAYER METAL4 ;
RECT 238.805 0.0 242.805 103.4 ;
LAYER METAL4 ;
RECT 227.185 0.0 231.185 103.4 ;
LAYER METAL4 ;
RECT 215.565 0.0 219.565 103.4 ;
LAYER METAL4 ;
RECT 203.945 0.0 207.945 103.4 ;
LAYER METAL4 ;
RECT 192.325 0.0 196.325 103.4 ;
LAYER METAL4 ;
RECT 180.705 0.0 184.705 103.4 ;
LAYER METAL4 ;
RECT 169.085 0.0 173.085 103.4 ;
LAYER METAL4 ;
RECT 157.465 0.0 161.465 103.4 ;
LAYER METAL4 ;
RECT 145.845 0.0 149.845 103.4 ;
LAYER METAL4 ;
RECT 134.225 0.0 138.225 103.4 ;
LAYER METAL4 ;
RECT 122.605 0.0 126.605 103.4 ;
LAYER METAL4 ;
RECT 110.985 0.0 114.985 103.4 ;
LAYER METAL4 ;
RECT 99.365 0.0 103.365 103.4 ;
LAYER METAL4 ;
RECT 87.745 0.0 91.745 103.4 ;
LAYER METAL4 ;
RECT 76.125 0.0 80.125 103.4 ;
LAYER METAL4 ;
RECT 64.505 0.0 68.505 103.4 ;
LAYER METAL4 ;
RECT 52.885 0.0 56.885 103.4 ;
LAYER METAL4 ;
RECT 41.265 0.0 45.265 103.4 ;
LAYER METAL4 ;
RECT 29.645 0.0 33.645 103.4 ;
LAYER METAL4 ;
RECT 18.025 0.0 22.025 103.4 ;
LAYER METAL4 ;
RECT 6.405 0.0 10.405 103.4 ;
LAYER METAL4 ;
RECT 387.475 0.0 391.475 103.4 ;
LAYER METAL4 ;
RECT 399.095 0.0 403.095 103.4 ;
LAYER METAL4 ;
RECT 410.715 0.0 414.715 103.4 ;
LAYER METAL4 ;
RECT 422.335 0.0 426.335 103.4 ;
LAYER METAL4 ;
RECT 433.955 0.0 437.955 103.4 ;
LAYER METAL4 ;
RECT 445.575 0.0 449.575 103.4 ;
LAYER METAL4 ;
RECT 457.195 0.0 461.195 103.4 ;
LAYER METAL4 ;
RECT 468.815 0.0 472.815 103.4 ;
LAYER METAL4 ;
RECT 480.435 0.0 484.435 103.4 ;
LAYER METAL4 ;
RECT 492.055 0.0 496.055 103.4 ;
LAYER METAL4 ;
RECT 503.675 0.0 507.675 103.4 ;
LAYER METAL4 ;
RECT 515.295 0.0 519.295 103.4 ;
LAYER METAL4 ;
RECT 526.915 0.0 530.915 103.4 ;
LAYER METAL4 ;
RECT 538.535 0.0 542.535 103.4 ;
LAYER METAL4 ;
RECT 550.155 0.0 554.155 103.4 ;
LAYER METAL4 ;
RECT 561.775 0.0 565.775 103.4 ;
LAYER METAL4 ;
RECT 573.395 0.0 577.395 103.4 ;
LAYER METAL4 ;
RECT 585.015 0.0 589.015 103.4 ;
LAYER METAL4 ;
RECT 596.635 0.0 600.635 103.4 ;
LAYER METAL4 ;
RECT 608.255 0.0 612.255 103.4 ;
LAYER METAL4 ;
RECT 619.875 0.0 623.875 103.4 ;
LAYER METAL4 ;
RECT 631.495 0.0 635.495 103.4 ;
LAYER METAL4 ;
RECT 643.115 0.0 647.115 103.4 ;
LAYER METAL4 ;
RECT 654.735 0.0 658.735 103.4 ;
END
END VDD

OBS
LAYER VIA12 ;
RECT  0.000 0.000 665.140 103.400 ;
LAYER VIA23 ;
RECT  0.000 0.000 665.140 103.400 ;
LAYER VIA34 ;
RECT  0.000 0.000 665.140 103.400 ;
LAYER METAL1 ;
POLYGON 0.000 0.000 18.495 0.000 18.495 0.870 20.025 0.870 20.025 0.000
 41.735 0.000 41.735 0.870 43.265 0.870 43.265 0.000 64.975 0.000
 64.975 0.870 66.505 0.870 66.505 0.000 88.215 0.000 88.215 0.870
 89.745 0.870 89.745 0.000 111.455 0.000 111.455 0.870 112.985 0.870
 112.985 0.000 134.695 0.000 134.695 0.870 136.225 0.870 136.225 0.000
 157.935 0.000 157.935 0.870 159.465 0.870 159.465 0.000 181.175 0.000
 181.175 0.870 182.705 0.870 182.705 0.000 204.415 0.000 204.415 0.870
 205.945 0.870 205.945 0.000 227.655 0.000 227.655 0.870 229.185 0.870
 229.185 0.000 250.895 0.000 250.895 0.870 252.425 0.870 252.425 0.000
 274.135 0.000 274.135 0.870 275.665 0.870 275.665 0.000 296.875 0.000
 296.875 1.300 297.835 1.300 297.835 0.000 306.490 0.000 306.490 1.300
 307.450 1.300 307.450 0.000 323.220 0.000 323.220 0.870 325.245 0.870
 325.245 0.000 328.980 0.000 328.980 0.870 331.005 0.870 331.005 0.000
 334.505 0.000 334.505 0.870 336.615 0.870 336.615 0.000 342.445 0.000
 342.445 0.870 344.555 0.870 344.555 0.000 350.385 0.000 350.385 0.870
 352.495 0.870 352.495 0.000 361.155 0.000 361.155 0.870 362.865 0.870
 362.865 0.000 366.005 0.000 366.005 0.870 367.715 0.870 367.715 0.000
 389.475 0.000 389.475 0.870 391.005 0.870 391.005 0.000 412.715 0.000
 412.715 0.870 414.245 0.870 414.245 0.000 435.955 0.000 435.955 0.870
 437.485 0.870 437.485 0.000 459.195 0.000 459.195 0.870 460.725 0.870
 460.725 0.000 482.435 0.000 482.435 0.870 483.965 0.870 483.965 0.000
 505.675 0.000 505.675 0.870 507.205 0.870 507.205 0.000 528.915 0.000
 528.915 0.870 530.445 0.870 530.445 0.000 552.155 0.000 552.155 0.870
 553.685 0.870 553.685 0.000 575.395 0.000 575.395 0.870 576.925 0.870
 576.925 0.000 598.635 0.000 598.635 0.870 600.165 0.870 600.165 0.000
 621.875 0.000 621.875 0.870 623.405 0.870 623.405 0.000 645.115 0.000
 645.115 0.870 646.645 0.870 646.645 0.000 665.140 0.000 665.140 103.400 656.465 103.400 656.465 102.530 654.935 102.530 654.935 103.400
 633.225 103.400 633.225 102.530 631.695 102.530 631.695 103.400 609.985 103.400
 609.985 102.530 608.455 102.530 608.455 103.400 586.745 103.400 586.745 102.530
 585.215 102.530 585.215 103.400 563.505 103.400 563.505 102.530 561.975 102.530
 561.975 103.400 540.265 103.400 540.265 102.530 538.735 102.530 538.735 103.400
 517.025 103.400 517.025 102.530 515.495 102.530 515.495 103.400 493.785 103.400
 493.785 102.530 492.255 102.530 492.255 103.400 470.545 103.400 470.545 102.530
 469.015 102.530 469.015 103.400 447.305 103.400 447.305 102.530 445.775 102.530
 445.775 103.400 424.065 103.400 424.065 102.530 422.535 102.530 422.535 103.400
 400.825 103.400 400.825 102.530 399.295 102.530 399.295 103.400 369.900 103.400
 369.900 102.100 368.940 102.100 368.940 103.400 360.495 103.400 360.495 102.100
 359.535 102.100 359.535 103.400 341.920 103.400 341.920 102.530 339.895 102.530
 339.895 103.400 336.160 103.400 336.160 102.530 334.135 102.530 334.135 103.400
 330.635 103.400 330.635 102.530 328.525 102.530 328.525 103.400 322.695 103.400
 322.695 102.530 320.585 102.530 320.585 103.400 314.755 103.400 314.755 102.530
 312.645 102.530 312.645 103.400 303.985 103.400 303.985 102.530 302.275 102.530
 302.275 103.400 299.135 103.400 299.135 102.530 297.425 102.530 297.425 103.400
 265.845 103.400 265.845 102.530 264.315 102.530 264.315 103.400 242.605 103.400
 242.605 102.530 241.075 102.530 241.075 103.400 219.365 103.400 219.365 102.530
 217.835 102.530 217.835 103.400 196.125 103.400 196.125 102.530 194.595 102.530
 194.595 103.400 172.885 103.400 172.885 102.530 171.355 102.530 171.355 103.400
 149.645 103.400 149.645 102.530 148.115 102.530 148.115 103.400 126.405 103.400
 126.405 102.530 124.875 102.530 124.875 103.400 103.165 103.400 103.165 102.530
 101.635 102.530 101.635 103.400 79.925 103.400 79.925 102.530 78.395 102.530
 78.395 103.400 56.685 103.400 56.685 102.530 55.155 102.530 55.155 103.400
 33.445 103.400 33.445 102.530 31.915 102.530 31.915 103.400 10.205 103.400
 10.205 102.530 8.675 102.530 8.675 103.400 0.000 103.400 ;
LAYER METAL2 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 334.855 0.000 334.855 0.920 336.665 0.920 336.665 0.000 342.795 0.000
 342.795 0.920 344.605 0.920 344.605 0.000 350.735 0.000 350.735 0.920
 352.545 0.920 352.545 0.000 361.105 0.000 361.105 0.920 362.915 0.920
 362.915 0.000 365.955 0.000 365.955 0.920 367.765 0.920 367.765 0.000
 389.425 0.000 389.425 0.920 391.055 0.920 391.055 0.000 412.665 0.000
 412.665 0.920 414.295 0.920 414.295 0.000 435.905 0.000 435.905 0.920
 437.535 0.920 437.535 0.000 459.145 0.000 459.145 0.920 460.775 0.920
 460.775 0.000 482.385 0.000 482.385 0.920 484.015 0.920 484.015 0.000
 505.625 0.000 505.625 0.920 507.255 0.920 507.255 0.000 528.865 0.000
 528.865 0.920 530.495 0.920 530.495 0.000 552.105 0.000 552.105 0.920
 553.735 0.920 553.735 0.000 575.345 0.000 575.345 0.920 576.975 0.920
 576.975 0.000 598.585 0.000 598.585 0.920 600.215 0.920 600.215 0.000
 621.825 0.000 621.825 0.920 623.455 0.920 623.455 0.000 645.065 0.000
 645.065 0.920 646.695 0.920 646.695 0.000 665.140 0.000 665.140 103.400 656.515 103.400 656.515 102.480 654.885 102.480 654.885 103.400
 633.275 103.400 633.275 102.480 631.645 102.480 631.645 103.400 610.035 103.400
 610.035 102.480 608.405 102.480 608.405 103.400 586.795 103.400 586.795 102.480
 585.165 102.480 585.165 103.400 563.555 103.400 563.555 102.480 561.925 102.480
 561.925 103.400 540.315 103.400 540.315 102.480 538.685 102.480 538.685 103.400
 517.075 103.400 517.075 102.480 515.445 102.480 515.445 103.400 493.835 103.400
 493.835 102.480 492.205 102.480 492.205 103.400 470.595 103.400 470.595 102.480
 468.965 102.480 468.965 103.400 447.355 103.400 447.355 102.480 445.725 102.480
 445.725 103.400 424.115 103.400 424.115 102.480 422.485 102.480 422.485 103.400
 400.875 103.400 400.875 102.480 399.245 102.480 399.245 103.400 369.950 103.400
 369.950 102.050 368.890 102.050 368.890 103.400 360.545 103.400 360.545 102.050
 359.485 102.050 359.485 103.400 341.655 103.400 341.655 102.480 339.845 102.480
 339.845 103.400 335.895 103.400 335.895 102.480 334.085 102.480 334.085 103.400
 330.285 103.400 330.285 102.480 328.475 102.480 328.475 103.400 322.345 103.400
 322.345 102.480 320.535 102.480 320.535 103.400 314.405 103.400 314.405 102.480
 312.595 102.480 312.595 103.400 304.035 103.400 304.035 102.480 302.225 102.480
 302.225 103.400 299.185 103.400 299.185 102.480 297.375 102.480 297.375 103.400
 265.895 103.400 265.895 102.480 264.265 102.480 264.265 103.400 242.655 103.400
 242.655 102.480 241.025 102.480 241.025 103.400 219.415 103.400 219.415 102.480
 217.785 102.480 217.785 103.400 196.175 103.400 196.175 102.480 194.545 102.480
 194.545 103.400 172.935 103.400 172.935 102.480 171.305 102.480 171.305 103.400
 149.695 103.400 149.695 102.480 148.065 102.480 148.065 103.400 126.455 103.400
 126.455 102.480 124.825 102.480 124.825 103.400 103.215 103.400 103.215 102.480
 101.585 102.480 101.585 103.400 79.975 103.400 79.975 102.480 78.345 102.480
 78.345 103.400 56.735 103.400 56.735 102.480 55.105 102.480 55.105 103.400
 33.495 103.400 33.495 102.480 31.865 102.480 31.865 103.400 10.255 103.400
 10.255 102.480 8.625 102.480 8.625 103.400 0.000 103.400 ;
LAYER METAL3 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 334.855 0.000 334.855 0.920 336.665 0.920 336.665 0.000 342.795 0.000
 342.795 0.920 344.605 0.920 344.605 0.000 350.735 0.000 350.735 0.920
 352.545 0.920 352.545 0.000 361.105 0.000 361.105 0.920 362.915 0.920
 362.915 0.000 365.955 0.000 365.955 0.920 367.765 0.920 367.765 0.000
 389.425 0.000 389.425 0.920 391.055 0.920 391.055 0.000 412.665 0.000
 412.665 0.920 414.295 0.920 414.295 0.000 435.905 0.000 435.905 0.920
 437.535 0.920 437.535 0.000 459.145 0.000 459.145 0.920 460.775 0.920
 460.775 0.000 482.385 0.000 482.385 0.920 484.015 0.920 484.015 0.000
 505.625 0.000 505.625 0.920 507.255 0.920 507.255 0.000 528.865 0.000
 528.865 0.920 530.495 0.920 530.495 0.000 552.105 0.000 552.105 0.920
 553.735 0.920 553.735 0.000 575.345 0.000 575.345 0.920 576.975 0.920
 576.975 0.000 598.585 0.000 598.585 0.920 600.215 0.920 600.215 0.000
 621.825 0.000 621.825 0.920 623.455 0.920 623.455 0.000 645.065 0.000
 645.065 0.920 646.695 0.920 646.695 0.000 665.140 0.000 665.140 103.400 656.515 103.400 656.515 102.480 654.885 102.480 654.885 103.400
 633.275 103.400 633.275 102.480 631.645 102.480 631.645 103.400 610.035 103.400
 610.035 102.480 608.405 102.480 608.405 103.400 586.795 103.400 586.795 102.480
 585.165 102.480 585.165 103.400 563.555 103.400 563.555 102.480 561.925 102.480
 561.925 103.400 540.315 103.400 540.315 102.480 538.685 102.480 538.685 103.400
 517.075 103.400 517.075 102.480 515.445 102.480 515.445 103.400 493.835 103.400
 493.835 102.480 492.205 102.480 492.205 103.400 470.595 103.400 470.595 102.480
 468.965 102.480 468.965 103.400 447.355 103.400 447.355 102.480 445.725 102.480
 445.725 103.400 424.115 103.400 424.115 102.480 422.485 102.480 422.485 103.400
 400.875 103.400 400.875 102.480 399.245 102.480 399.245 103.400 369.950 103.400
 369.950 102.050 368.890 102.050 368.890 103.400 360.545 103.400 360.545 102.050
 359.485 102.050 359.485 103.400 341.655 103.400 341.655 102.480 339.845 102.480
 339.845 103.400 335.895 103.400 335.895 102.480 334.085 102.480 334.085 103.400
 330.285 103.400 330.285 102.480 328.475 102.480 328.475 103.400 322.345 103.400
 322.345 102.480 320.535 102.480 320.535 103.400 314.405 103.400 314.405 102.480
 312.595 102.480 312.595 103.400 304.035 103.400 304.035 102.480 302.225 102.480
 302.225 103.400 299.185 103.400 299.185 102.480 297.375 102.480 297.375 103.400
 265.895 103.400 265.895 102.480 264.265 102.480 264.265 103.400 242.655 103.400
 242.655 102.480 241.025 102.480 241.025 103.400 219.415 103.400 219.415 102.480
 217.785 102.480 217.785 103.400 196.175 103.400 196.175 102.480 194.545 102.480
 194.545 103.400 172.935 103.400 172.935 102.480 171.305 102.480 171.305 103.400
 149.695 103.400 149.695 102.480 148.065 102.480 148.065 103.400 126.455 103.400
 126.455 102.480 124.825 102.480 124.825 103.400 103.215 103.400 103.215 102.480
 101.585 102.480 101.585 103.400 79.975 103.400 79.975 102.480 78.345 102.480
 78.345 103.400 56.735 103.400 56.735 102.480 55.105 102.480 55.105 103.400
 33.495 103.400 33.495 102.480 31.865 102.480 31.865 103.400 10.255 103.400
 10.255 102.480 8.625 102.480 8.625 103.400 0.000 103.400 ;
END
END RAM128
END LIBRARY
