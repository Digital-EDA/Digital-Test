************************************************************************
* auCdl Netlist:
*
* Library Name:  SMIC_MEMORY
* Top Cell Name: FRAM512
* Version:  V0.2
* View Name:     schematic
* Netlisted on:  Wed May 31 22:22:18 CST 2023
************************************************************************
*.BIPOLAR
*.RESI = 2000
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM


************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELLDBL
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELLDBL BB VDD VSS
MM4 BB VSS VSS VSS N18 W=220.00N L=225.00N M=1
MM1 VSS VSS VSS VSS N18 W=705.00N L=180.00N M=1
MM7 VSS VSS VSS VSS N18 W=220.00N L=225.00N M=1
MM6 VDD VDD VDD VDD P18 W=220.000N L=200.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL_EDGE256
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL_EDGE256 DBL VDD VSS
XI0 DBL VDD VSS FRAM512_BITCELLDBL
XI1 DBL VDD VSS FRAM512_BITCELLDBL
XI2 DBL VDD VSS FRAM512_BITCELLDBL
XI3 DBL VDD VSS FRAM512_BITCELLDBL
XI4 DBL VDD VSS FRAM512_BITCELLDBL
XI5 DBL VDD VSS FRAM512_BITCELLDBL
XI6 DBL VDD VSS FRAM512_BITCELLDBL
XI7 DBL VDD VSS FRAM512_BITCELLDBL
XI8 DBL VDD VSS FRAM512_BITCELLDBL
XI9 DBL VDD VSS FRAM512_BITCELLDBL
XI10 DBL VDD VSS FRAM512_BITCELLDBL
XI11 DBL VDD VSS FRAM512_BITCELLDBL
XI12 DBL VDD VSS FRAM512_BITCELLDBL
XI13 DBL VDD VSS FRAM512_BITCELLDBL
XI14 DBL VDD VSS FRAM512_BITCELLDBL
XI15 DBL VDD VSS FRAM512_BITCELLDBL
XI16 DBL VDD VSS FRAM512_BITCELLDBL
XI17 DBL VDD VSS FRAM512_BITCELLDBL
XI18 DBL VDD VSS FRAM512_BITCELLDBL
XI19 DBL VDD VSS FRAM512_BITCELLDBL
XI20 DBL VDD VSS FRAM512_BITCELLDBL
XI21 DBL VDD VSS FRAM512_BITCELLDBL
XI22 DBL VDD VSS FRAM512_BITCELLDBL
XI23 DBL VDD VSS FRAM512_BITCELLDBL
XI24 DBL VDD VSS FRAM512_BITCELLDBL
XI25 DBL VDD VSS FRAM512_BITCELLDBL
XI26 DBL VDD VSS FRAM512_BITCELLDBL
XI27 DBL VDD VSS FRAM512_BITCELLDBL
XI28 DBL VDD VSS FRAM512_BITCELLDBL
XI29 DBL VDD VSS FRAM512_BITCELLDBL
XI30 DBL VDD VSS FRAM512_BITCELLDBL
XI31 DBL VDD VSS FRAM512_BITCELLDBL
XI32 DBL VDD VSS FRAM512_BITCELLDBL
XI33 DBL VDD VSS FRAM512_BITCELLDBL
XI34 DBL VDD VSS FRAM512_BITCELLDBL
XI35 DBL VDD VSS FRAM512_BITCELLDBL
XI36 DBL VDD VSS FRAM512_BITCELLDBL
XI37 DBL VDD VSS FRAM512_BITCELLDBL
XI38 DBL VDD VSS FRAM512_BITCELLDBL
XI39 DBL VDD VSS FRAM512_BITCELLDBL
XI40 DBL VDD VSS FRAM512_BITCELLDBL
XI41 DBL VDD VSS FRAM512_BITCELLDBL
XI42 DBL VDD VSS FRAM512_BITCELLDBL
XI43 DBL VDD VSS FRAM512_BITCELLDBL
XI44 DBL VDD VSS FRAM512_BITCELLDBL
XI45 DBL VDD VSS FRAM512_BITCELLDBL
XI46 DBL VDD VSS FRAM512_BITCELLDBL
XI47 DBL VDD VSS FRAM512_BITCELLDBL
XI48 DBL VDD VSS FRAM512_BITCELLDBL
XI49 DBL VDD VSS FRAM512_BITCELLDBL
XI50 DBL VDD VSS FRAM512_BITCELLDBL
XI51 DBL VDD VSS FRAM512_BITCELLDBL
XI52 DBL VDD VSS FRAM512_BITCELLDBL
XI53 DBL VDD VSS FRAM512_BITCELLDBL
XI54 DBL VDD VSS FRAM512_BITCELLDBL
XI55 DBL VDD VSS FRAM512_BITCELLDBL
XI56 DBL VDD VSS FRAM512_BITCELLDBL
XI57 DBL VDD VSS FRAM512_BITCELLDBL
XI58 DBL VDD VSS FRAM512_BITCELLDBL
XI59 DBL VDD VSS FRAM512_BITCELLDBL
XI60 DBL VDD VSS FRAM512_BITCELLDBL
XI61 DBL VDD VSS FRAM512_BITCELLDBL
XI62 DBL VDD VSS FRAM512_BITCELLDBL
XI63 DBL VDD VSS FRAM512_BITCELLDBL
XI64 DBL VDD VSS FRAM512_BITCELLDBL
XI65 DBL VDD VSS FRAM512_BITCELLDBL
XI66 DBL VDD VSS FRAM512_BITCELLDBL
XI67 DBL VDD VSS FRAM512_BITCELLDBL
XI68 DBL VDD VSS FRAM512_BITCELLDBL
XI69 DBL VDD VSS FRAM512_BITCELLDBL
XI70 DBL VDD VSS FRAM512_BITCELLDBL
XI71 DBL VDD VSS FRAM512_BITCELLDBL
XI72 DBL VDD VSS FRAM512_BITCELLDBL
XI73 DBL VDD VSS FRAM512_BITCELLDBL
XI74 DBL VDD VSS FRAM512_BITCELLDBL
XI75 DBL VDD VSS FRAM512_BITCELLDBL
XI76 DBL VDD VSS FRAM512_BITCELLDBL
XI77 DBL VDD VSS FRAM512_BITCELLDBL
XI78 DBL VDD VSS FRAM512_BITCELLDBL
XI79 DBL VDD VSS FRAM512_BITCELLDBL
XI80 DBL VDD VSS FRAM512_BITCELLDBL
XI81 DBL VDD VSS FRAM512_BITCELLDBL
XI82 DBL VDD VSS FRAM512_BITCELLDBL
XI83 DBL VDD VSS FRAM512_BITCELLDBL
XI84 DBL VDD VSS FRAM512_BITCELLDBL
XI85 DBL VDD VSS FRAM512_BITCELLDBL
XI86 DBL VDD VSS FRAM512_BITCELLDBL
XI87 DBL VDD VSS FRAM512_BITCELLDBL
XI88 DBL VDD VSS FRAM512_BITCELLDBL
XI89 DBL VDD VSS FRAM512_BITCELLDBL
XI90 DBL VDD VSS FRAM512_BITCELLDBL
XI91 DBL VDD VSS FRAM512_BITCELLDBL
XI92 DBL VDD VSS FRAM512_BITCELLDBL
XI93 DBL VDD VSS FRAM512_BITCELLDBL
XI94 DBL VDD VSS FRAM512_BITCELLDBL
XI95 DBL VDD VSS FRAM512_BITCELLDBL
XI96 DBL VDD VSS FRAM512_BITCELLDBL
XI97 DBL VDD VSS FRAM512_BITCELLDBL
XI98 DBL VDD VSS FRAM512_BITCELLDBL
XI99 DBL VDD VSS FRAM512_BITCELLDBL
XI100 DBL VDD VSS FRAM512_BITCELLDBL
XI101 DBL VDD VSS FRAM512_BITCELLDBL
XI102 DBL VDD VSS FRAM512_BITCELLDBL
XI103 DBL VDD VSS FRAM512_BITCELLDBL
XI104 DBL VDD VSS FRAM512_BITCELLDBL
XI105 DBL VDD VSS FRAM512_BITCELLDBL
XI106 DBL VDD VSS FRAM512_BITCELLDBL
XI107 DBL VDD VSS FRAM512_BITCELLDBL
XI108 DBL VDD VSS FRAM512_BITCELLDBL
XI109 DBL VDD VSS FRAM512_BITCELLDBL
XI110 DBL VDD VSS FRAM512_BITCELLDBL
XI111 DBL VDD VSS FRAM512_BITCELLDBL
XI112 DBL VDD VSS FRAM512_BITCELLDBL
XI113 DBL VDD VSS FRAM512_BITCELLDBL
XI114 DBL VDD VSS FRAM512_BITCELLDBL
XI115 DBL VDD VSS FRAM512_BITCELLDBL
XI116 DBL VDD VSS FRAM512_BITCELLDBL
XI117 DBL VDD VSS FRAM512_BITCELLDBL
XI118 DBL VDD VSS FRAM512_BITCELLDBL
XI119 DBL VDD VSS FRAM512_BITCELLDBL
XI120 DBL VDD VSS FRAM512_BITCELLDBL
XI121 DBL VDD VSS FRAM512_BITCELLDBL
XI122 DBL VDD VSS FRAM512_BITCELLDBL
XI123 DBL VDD VSS FRAM512_BITCELLDBL
XI124 DBL VDD VSS FRAM512_BITCELLDBL
XI125 DBL VDD VSS FRAM512_BITCELLDBL
XI126 DBL VDD VSS FRAM512_BITCELLDBL
XI127 DBL VDD VSS FRAM512_BITCELLDBL
XI128 DBL VDD VSS FRAM512_BITCELLDBL
XI129 DBL VDD VSS FRAM512_BITCELLDBL
XI130 DBL VDD VSS FRAM512_BITCELLDBL
XI131 DBL VDD VSS FRAM512_BITCELLDBL
XI132 DBL VDD VSS FRAM512_BITCELLDBL
XI133 DBL VDD VSS FRAM512_BITCELLDBL
XI134 DBL VDD VSS FRAM512_BITCELLDBL
XI135 DBL VDD VSS FRAM512_BITCELLDBL
XI136 DBL VDD VSS FRAM512_BITCELLDBL
XI137 DBL VDD VSS FRAM512_BITCELLDBL
XI138 DBL VDD VSS FRAM512_BITCELLDBL
XI139 DBL VDD VSS FRAM512_BITCELLDBL
XI140 DBL VDD VSS FRAM512_BITCELLDBL
XI141 DBL VDD VSS FRAM512_BITCELLDBL
XI142 DBL VDD VSS FRAM512_BITCELLDBL
XI143 DBL VDD VSS FRAM512_BITCELLDBL
XI144 DBL VDD VSS FRAM512_BITCELLDBL
XI145 DBL VDD VSS FRAM512_BITCELLDBL
XI146 DBL VDD VSS FRAM512_BITCELLDBL
XI147 DBL VDD VSS FRAM512_BITCELLDBL
XI148 DBL VDD VSS FRAM512_BITCELLDBL
XI149 DBL VDD VSS FRAM512_BITCELLDBL
XI150 DBL VDD VSS FRAM512_BITCELLDBL
XI151 DBL VDD VSS FRAM512_BITCELLDBL
XI152 DBL VDD VSS FRAM512_BITCELLDBL
XI153 DBL VDD VSS FRAM512_BITCELLDBL
XI154 DBL VDD VSS FRAM512_BITCELLDBL
XI155 DBL VDD VSS FRAM512_BITCELLDBL
XI156 DBL VDD VSS FRAM512_BITCELLDBL
XI157 DBL VDD VSS FRAM512_BITCELLDBL
XI158 DBL VDD VSS FRAM512_BITCELLDBL
XI159 DBL VDD VSS FRAM512_BITCELLDBL
XI160 DBL VDD VSS FRAM512_BITCELLDBL
XI161 DBL VDD VSS FRAM512_BITCELLDBL
XI162 DBL VDD VSS FRAM512_BITCELLDBL
XI163 DBL VDD VSS FRAM512_BITCELLDBL
XI164 DBL VDD VSS FRAM512_BITCELLDBL
XI165 DBL VDD VSS FRAM512_BITCELLDBL
XI166 DBL VDD VSS FRAM512_BITCELLDBL
XI167 DBL VDD VSS FRAM512_BITCELLDBL
XI168 DBL VDD VSS FRAM512_BITCELLDBL
XI169 DBL VDD VSS FRAM512_BITCELLDBL
XI170 DBL VDD VSS FRAM512_BITCELLDBL
XI171 DBL VDD VSS FRAM512_BITCELLDBL
XI172 DBL VDD VSS FRAM512_BITCELLDBL
XI173 DBL VDD VSS FRAM512_BITCELLDBL
XI174 DBL VDD VSS FRAM512_BITCELLDBL
XI175 DBL VDD VSS FRAM512_BITCELLDBL
XI176 DBL VDD VSS FRAM512_BITCELLDBL
XI177 DBL VDD VSS FRAM512_BITCELLDBL
XI178 DBL VDD VSS FRAM512_BITCELLDBL
XI179 DBL VDD VSS FRAM512_BITCELLDBL
XI180 DBL VDD VSS FRAM512_BITCELLDBL
XI181 DBL VDD VSS FRAM512_BITCELLDBL
XI182 DBL VDD VSS FRAM512_BITCELLDBL
XI183 DBL VDD VSS FRAM512_BITCELLDBL
XI184 DBL VDD VSS FRAM512_BITCELLDBL
XI185 DBL VDD VSS FRAM512_BITCELLDBL
XI186 DBL VDD VSS FRAM512_BITCELLDBL
XI187 DBL VDD VSS FRAM512_BITCELLDBL
XI188 DBL VDD VSS FRAM512_BITCELLDBL
XI189 DBL VDD VSS FRAM512_BITCELLDBL
XI190 DBL VDD VSS FRAM512_BITCELLDBL
XI191 DBL VDD VSS FRAM512_BITCELLDBL
XI192 DBL VDD VSS FRAM512_BITCELLDBL
XI193 DBL VDD VSS FRAM512_BITCELLDBL
XI194 DBL VDD VSS FRAM512_BITCELLDBL
XI195 DBL VDD VSS FRAM512_BITCELLDBL
XI196 DBL VDD VSS FRAM512_BITCELLDBL
XI197 DBL VDD VSS FRAM512_BITCELLDBL
XI198 DBL VDD VSS FRAM512_BITCELLDBL
XI199 DBL VDD VSS FRAM512_BITCELLDBL
XI200 DBL VDD VSS FRAM512_BITCELLDBL
XI201 DBL VDD VSS FRAM512_BITCELLDBL
XI202 DBL VDD VSS FRAM512_BITCELLDBL
XI203 DBL VDD VSS FRAM512_BITCELLDBL
XI204 DBL VDD VSS FRAM512_BITCELLDBL
XI205 DBL VDD VSS FRAM512_BITCELLDBL
XI206 DBL VDD VSS FRAM512_BITCELLDBL
XI207 DBL VDD VSS FRAM512_BITCELLDBL
XI208 DBL VDD VSS FRAM512_BITCELLDBL
XI209 DBL VDD VSS FRAM512_BITCELLDBL
XI210 DBL VDD VSS FRAM512_BITCELLDBL
XI211 DBL VDD VSS FRAM512_BITCELLDBL
XI212 DBL VDD VSS FRAM512_BITCELLDBL
XI213 DBL VDD VSS FRAM512_BITCELLDBL
XI214 DBL VDD VSS FRAM512_BITCELLDBL
XI215 DBL VDD VSS FRAM512_BITCELLDBL
XI216 DBL VDD VSS FRAM512_BITCELLDBL
XI217 DBL VDD VSS FRAM512_BITCELLDBL
XI218 DBL VDD VSS FRAM512_BITCELLDBL
XI219 DBL VDD VSS FRAM512_BITCELLDBL
XI220 DBL VDD VSS FRAM512_BITCELLDBL
XI221 DBL VDD VSS FRAM512_BITCELLDBL
XI222 DBL VDD VSS FRAM512_BITCELLDBL
XI223 DBL VDD VSS FRAM512_BITCELLDBL
XI224 DBL VDD VSS FRAM512_BITCELLDBL
XI225 DBL VDD VSS FRAM512_BITCELLDBL
XI226 DBL VDD VSS FRAM512_BITCELLDBL
XI227 DBL VDD VSS FRAM512_BITCELLDBL
XI228 DBL VDD VSS FRAM512_BITCELLDBL
XI229 DBL VDD VSS FRAM512_BITCELLDBL
XI230 DBL VDD VSS FRAM512_BITCELLDBL
XI231 DBL VDD VSS FRAM512_BITCELLDBL
XI232 DBL VDD VSS FRAM512_BITCELLDBL
XI233 DBL VDD VSS FRAM512_BITCELLDBL
XI234 DBL VDD VSS FRAM512_BITCELLDBL
XI235 DBL VDD VSS FRAM512_BITCELLDBL
XI236 DBL VDD VSS FRAM512_BITCELLDBL
XI237 DBL VDD VSS FRAM512_BITCELLDBL
XI238 DBL VDD VSS FRAM512_BITCELLDBL
XI239 DBL VDD VSS FRAM512_BITCELLDBL
XI240 DBL VDD VSS FRAM512_BITCELLDBL
XI241 DBL VDD VSS FRAM512_BITCELLDBL
XI242 DBL VDD VSS FRAM512_BITCELLDBL
XI243 DBL VDD VSS FRAM512_BITCELLDBL
XI244 DBL VDD VSS FRAM512_BITCELLDBL
XI245 DBL VDD VSS FRAM512_BITCELLDBL
XI246 DBL VDD VSS FRAM512_BITCELLDBL
XI247 DBL VDD VSS FRAM512_BITCELLDBL
XI248 DBL VDD VSS FRAM512_BITCELLDBL
XI249 DBL VDD VSS FRAM512_BITCELLDBL
XI250 DBL VDD VSS FRAM512_BITCELLDBL
XI251 DBL VDD VSS FRAM512_BITCELLDBL
XI252 DBL VDD VSS FRAM512_BITCELLDBL
XI253 DBL VDD VSS FRAM512_BITCELLDBL
XI254 DBL VDD VSS FRAM512_BITCELLDBL
XI255 DBL VDD VSS FRAM512_BITCELLDBL
XI256 NET12 VDD VSS FRAM512_BITCELLDBL
XI257 NET12 VDD VSS FRAM512_BITCELLDBL
XI258 NET18 VDD VSS FRAM512_BITCELLDBL
XI259 DBL VDD VSS FRAM512_BITCELLDBL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELLDUM
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELLDUM VSS WLA
MM4 VSS WLA VSS VSS N18 W=220.00N L=225.00N M=1
MM1 VSS VSS VSS VSS N18 W=705.00N L=180.00N M=1
MM7 VSS WLA VSS VSS N18 W=220.00N L=225.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_PCAP_DUMMY256
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_PCAP_DUMMY256 STWL[3] STWL[2] STWL[1] STWL[0] VSS WL[255] WL[254] WL[253] WL[252] WL[251]
+WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231]
+WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221]
+WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211]
+WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191]
+WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181]
+WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171]
+WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151]
+WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141]
+WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131]
+WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111]
+WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101]
+WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91]
+WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71]
+WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
XI0 VSS WL[255] FRAM512_BITCELLDUM
XI1 VSS WL[254] FRAM512_BITCELLDUM
XI2 VSS WL[253] FRAM512_BITCELLDUM
XI3 VSS WL[252] FRAM512_BITCELLDUM
XI4 VSS WL[251] FRAM512_BITCELLDUM
XI5 VSS WL[250] FRAM512_BITCELLDUM
XI6 VSS WL[249] FRAM512_BITCELLDUM
XI7 VSS WL[248] FRAM512_BITCELLDUM
XI8 VSS WL[247] FRAM512_BITCELLDUM
XI9 VSS WL[246] FRAM512_BITCELLDUM
XI10 VSS WL[245] FRAM512_BITCELLDUM
XI11 VSS WL[244] FRAM512_BITCELLDUM
XI12 VSS WL[243] FRAM512_BITCELLDUM
XI13 VSS WL[242] FRAM512_BITCELLDUM
XI14 VSS WL[241] FRAM512_BITCELLDUM
XI15 VSS WL[240] FRAM512_BITCELLDUM
XI16 VSS WL[239] FRAM512_BITCELLDUM
XI17 VSS WL[238] FRAM512_BITCELLDUM
XI18 VSS WL[237] FRAM512_BITCELLDUM
XI19 VSS WL[236] FRAM512_BITCELLDUM
XI20 VSS WL[235] FRAM512_BITCELLDUM
XI21 VSS WL[234] FRAM512_BITCELLDUM
XI22 VSS WL[233] FRAM512_BITCELLDUM
XI23 VSS WL[232] FRAM512_BITCELLDUM
XI24 VSS WL[231] FRAM512_BITCELLDUM
XI25 VSS WL[230] FRAM512_BITCELLDUM
XI26 VSS WL[229] FRAM512_BITCELLDUM
XI27 VSS WL[228] FRAM512_BITCELLDUM
XI28 VSS WL[227] FRAM512_BITCELLDUM
XI29 VSS WL[226] FRAM512_BITCELLDUM
XI30 VSS WL[225] FRAM512_BITCELLDUM
XI31 VSS WL[224] FRAM512_BITCELLDUM
XI32 VSS WL[223] FRAM512_BITCELLDUM
XI33 VSS WL[222] FRAM512_BITCELLDUM
XI34 VSS WL[221] FRAM512_BITCELLDUM
XI35 VSS WL[220] FRAM512_BITCELLDUM
XI36 VSS WL[219] FRAM512_BITCELLDUM
XI37 VSS WL[218] FRAM512_BITCELLDUM
XI38 VSS WL[217] FRAM512_BITCELLDUM
XI39 VSS WL[216] FRAM512_BITCELLDUM
XI40 VSS WL[215] FRAM512_BITCELLDUM
XI41 VSS WL[214] FRAM512_BITCELLDUM
XI42 VSS WL[213] FRAM512_BITCELLDUM
XI43 VSS WL[212] FRAM512_BITCELLDUM
XI44 VSS WL[211] FRAM512_BITCELLDUM
XI45 VSS WL[210] FRAM512_BITCELLDUM
XI46 VSS WL[209] FRAM512_BITCELLDUM
XI47 VSS WL[208] FRAM512_BITCELLDUM
XI48 VSS WL[207] FRAM512_BITCELLDUM
XI49 VSS WL[206] FRAM512_BITCELLDUM
XI50 VSS WL[205] FRAM512_BITCELLDUM
XI51 VSS WL[204] FRAM512_BITCELLDUM
XI52 VSS WL[203] FRAM512_BITCELLDUM
XI53 VSS WL[202] FRAM512_BITCELLDUM
XI54 VSS WL[201] FRAM512_BITCELLDUM
XI55 VSS WL[200] FRAM512_BITCELLDUM
XI56 VSS WL[199] FRAM512_BITCELLDUM
XI57 VSS WL[198] FRAM512_BITCELLDUM
XI58 VSS WL[197] FRAM512_BITCELLDUM
XI59 VSS WL[196] FRAM512_BITCELLDUM
XI60 VSS WL[195] FRAM512_BITCELLDUM
XI61 VSS WL[194] FRAM512_BITCELLDUM
XI62 VSS WL[193] FRAM512_BITCELLDUM
XI63 VSS WL[192] FRAM512_BITCELLDUM
XI64 VSS WL[191] FRAM512_BITCELLDUM
XI65 VSS WL[190] FRAM512_BITCELLDUM
XI66 VSS WL[189] FRAM512_BITCELLDUM
XI67 VSS WL[188] FRAM512_BITCELLDUM
XI68 VSS WL[187] FRAM512_BITCELLDUM
XI69 VSS WL[186] FRAM512_BITCELLDUM
XI70 VSS WL[185] FRAM512_BITCELLDUM
XI71 VSS WL[184] FRAM512_BITCELLDUM
XI72 VSS WL[183] FRAM512_BITCELLDUM
XI73 VSS WL[182] FRAM512_BITCELLDUM
XI74 VSS WL[181] FRAM512_BITCELLDUM
XI75 VSS WL[180] FRAM512_BITCELLDUM
XI76 VSS WL[179] FRAM512_BITCELLDUM
XI77 VSS WL[178] FRAM512_BITCELLDUM
XI78 VSS WL[177] FRAM512_BITCELLDUM
XI79 VSS WL[176] FRAM512_BITCELLDUM
XI80 VSS WL[175] FRAM512_BITCELLDUM
XI81 VSS WL[174] FRAM512_BITCELLDUM
XI82 VSS WL[173] FRAM512_BITCELLDUM
XI83 VSS WL[172] FRAM512_BITCELLDUM
XI84 VSS WL[171] FRAM512_BITCELLDUM
XI85 VSS WL[170] FRAM512_BITCELLDUM
XI86 VSS WL[169] FRAM512_BITCELLDUM
XI87 VSS WL[168] FRAM512_BITCELLDUM
XI88 VSS WL[167] FRAM512_BITCELLDUM
XI89 VSS WL[166] FRAM512_BITCELLDUM
XI90 VSS WL[165] FRAM512_BITCELLDUM
XI91 VSS WL[164] FRAM512_BITCELLDUM
XI92 VSS WL[163] FRAM512_BITCELLDUM
XI93 VSS WL[162] FRAM512_BITCELLDUM
XI94 VSS WL[161] FRAM512_BITCELLDUM
XI95 VSS WL[160] FRAM512_BITCELLDUM
XI96 VSS WL[159] FRAM512_BITCELLDUM
XI97 VSS WL[158] FRAM512_BITCELLDUM
XI98 VSS WL[157] FRAM512_BITCELLDUM
XI99 VSS WL[156] FRAM512_BITCELLDUM
XI100 VSS WL[155] FRAM512_BITCELLDUM
XI101 VSS WL[154] FRAM512_BITCELLDUM
XI102 VSS WL[153] FRAM512_BITCELLDUM
XI103 VSS WL[152] FRAM512_BITCELLDUM
XI104 VSS WL[151] FRAM512_BITCELLDUM
XI105 VSS WL[150] FRAM512_BITCELLDUM
XI106 VSS WL[149] FRAM512_BITCELLDUM
XI107 VSS WL[148] FRAM512_BITCELLDUM
XI108 VSS WL[147] FRAM512_BITCELLDUM
XI109 VSS WL[146] FRAM512_BITCELLDUM
XI110 VSS WL[145] FRAM512_BITCELLDUM
XI111 VSS WL[144] FRAM512_BITCELLDUM
XI112 VSS WL[143] FRAM512_BITCELLDUM
XI113 VSS WL[142] FRAM512_BITCELLDUM
XI114 VSS WL[141] FRAM512_BITCELLDUM
XI115 VSS WL[140] FRAM512_BITCELLDUM
XI116 VSS WL[139] FRAM512_BITCELLDUM
XI117 VSS WL[138] FRAM512_BITCELLDUM
XI118 VSS WL[137] FRAM512_BITCELLDUM
XI119 VSS WL[136] FRAM512_BITCELLDUM
XI120 VSS WL[135] FRAM512_BITCELLDUM
XI121 VSS WL[134] FRAM512_BITCELLDUM
XI122 VSS WL[133] FRAM512_BITCELLDUM
XI123 VSS WL[132] FRAM512_BITCELLDUM
XI124 VSS WL[131] FRAM512_BITCELLDUM
XI125 VSS WL[130] FRAM512_BITCELLDUM
XI126 VSS WL[129] FRAM512_BITCELLDUM
XI127 VSS WL[128] FRAM512_BITCELLDUM
XI128 VSS WL[127] FRAM512_BITCELLDUM
XI129 VSS WL[126] FRAM512_BITCELLDUM
XI130 VSS WL[125] FRAM512_BITCELLDUM
XI131 VSS WL[124] FRAM512_BITCELLDUM
XI132 VSS WL[123] FRAM512_BITCELLDUM
XI133 VSS WL[122] FRAM512_BITCELLDUM
XI134 VSS WL[121] FRAM512_BITCELLDUM
XI135 VSS WL[120] FRAM512_BITCELLDUM
XI136 VSS WL[119] FRAM512_BITCELLDUM
XI137 VSS WL[118] FRAM512_BITCELLDUM
XI138 VSS WL[117] FRAM512_BITCELLDUM
XI139 VSS WL[116] FRAM512_BITCELLDUM
XI140 VSS WL[115] FRAM512_BITCELLDUM
XI141 VSS WL[114] FRAM512_BITCELLDUM
XI142 VSS WL[113] FRAM512_BITCELLDUM
XI143 VSS WL[112] FRAM512_BITCELLDUM
XI144 VSS WL[111] FRAM512_BITCELLDUM
XI145 VSS WL[110] FRAM512_BITCELLDUM
XI146 VSS WL[109] FRAM512_BITCELLDUM
XI147 VSS WL[108] FRAM512_BITCELLDUM
XI148 VSS WL[107] FRAM512_BITCELLDUM
XI149 VSS WL[106] FRAM512_BITCELLDUM
XI150 VSS WL[105] FRAM512_BITCELLDUM
XI151 VSS WL[104] FRAM512_BITCELLDUM
XI152 VSS WL[103] FRAM512_BITCELLDUM
XI153 VSS WL[102] FRAM512_BITCELLDUM
XI154 VSS WL[101] FRAM512_BITCELLDUM
XI155 VSS WL[100] FRAM512_BITCELLDUM
XI156 VSS WL[99] FRAM512_BITCELLDUM
XI157 VSS WL[98] FRAM512_BITCELLDUM
XI158 VSS WL[97] FRAM512_BITCELLDUM
XI159 VSS WL[96] FRAM512_BITCELLDUM
XI160 VSS WL[95] FRAM512_BITCELLDUM
XI161 VSS WL[94] FRAM512_BITCELLDUM
XI162 VSS WL[93] FRAM512_BITCELLDUM
XI163 VSS WL[92] FRAM512_BITCELLDUM
XI164 VSS WL[91] FRAM512_BITCELLDUM
XI165 VSS WL[90] FRAM512_BITCELLDUM
XI166 VSS WL[89] FRAM512_BITCELLDUM
XI167 VSS WL[88] FRAM512_BITCELLDUM
XI168 VSS WL[87] FRAM512_BITCELLDUM
XI169 VSS WL[86] FRAM512_BITCELLDUM
XI170 VSS WL[85] FRAM512_BITCELLDUM
XI171 VSS WL[84] FRAM512_BITCELLDUM
XI172 VSS WL[83] FRAM512_BITCELLDUM
XI173 VSS WL[82] FRAM512_BITCELLDUM
XI174 VSS WL[81] FRAM512_BITCELLDUM
XI175 VSS WL[80] FRAM512_BITCELLDUM
XI176 VSS WL[79] FRAM512_BITCELLDUM
XI177 VSS WL[78] FRAM512_BITCELLDUM
XI178 VSS WL[77] FRAM512_BITCELLDUM
XI179 VSS WL[76] FRAM512_BITCELLDUM
XI180 VSS WL[75] FRAM512_BITCELLDUM
XI181 VSS WL[74] FRAM512_BITCELLDUM
XI182 VSS WL[73] FRAM512_BITCELLDUM
XI183 VSS WL[72] FRAM512_BITCELLDUM
XI184 VSS WL[71] FRAM512_BITCELLDUM
XI185 VSS WL[70] FRAM512_BITCELLDUM
XI186 VSS WL[69] FRAM512_BITCELLDUM
XI187 VSS WL[68] FRAM512_BITCELLDUM
XI188 VSS WL[67] FRAM512_BITCELLDUM
XI189 VSS WL[66] FRAM512_BITCELLDUM
XI190 VSS WL[65] FRAM512_BITCELLDUM
XI191 VSS WL[64] FRAM512_BITCELLDUM
XI192 VSS WL[63] FRAM512_BITCELLDUM
XI193 VSS WL[62] FRAM512_BITCELLDUM
XI194 VSS WL[61] FRAM512_BITCELLDUM
XI195 VSS WL[60] FRAM512_BITCELLDUM
XI196 VSS WL[59] FRAM512_BITCELLDUM
XI197 VSS WL[58] FRAM512_BITCELLDUM
XI198 VSS WL[57] FRAM512_BITCELLDUM
XI199 VSS WL[56] FRAM512_BITCELLDUM
XI200 VSS WL[55] FRAM512_BITCELLDUM
XI201 VSS WL[54] FRAM512_BITCELLDUM
XI202 VSS WL[53] FRAM512_BITCELLDUM
XI203 VSS WL[52] FRAM512_BITCELLDUM
XI204 VSS WL[51] FRAM512_BITCELLDUM
XI205 VSS WL[50] FRAM512_BITCELLDUM
XI206 VSS WL[49] FRAM512_BITCELLDUM
XI207 VSS WL[48] FRAM512_BITCELLDUM
XI208 VSS WL[47] FRAM512_BITCELLDUM
XI209 VSS WL[46] FRAM512_BITCELLDUM
XI210 VSS WL[45] FRAM512_BITCELLDUM
XI211 VSS WL[44] FRAM512_BITCELLDUM
XI212 VSS WL[43] FRAM512_BITCELLDUM
XI213 VSS WL[42] FRAM512_BITCELLDUM
XI214 VSS WL[41] FRAM512_BITCELLDUM
XI215 VSS WL[40] FRAM512_BITCELLDUM
XI216 VSS WL[39] FRAM512_BITCELLDUM
XI217 VSS WL[38] FRAM512_BITCELLDUM
XI218 VSS WL[37] FRAM512_BITCELLDUM
XI219 VSS WL[36] FRAM512_BITCELLDUM
XI220 VSS WL[35] FRAM512_BITCELLDUM
XI221 VSS WL[34] FRAM512_BITCELLDUM
XI222 VSS WL[33] FRAM512_BITCELLDUM
XI223 VSS WL[32] FRAM512_BITCELLDUM
XI224 VSS WL[31] FRAM512_BITCELLDUM
XI225 VSS WL[30] FRAM512_BITCELLDUM
XI226 VSS WL[29] FRAM512_BITCELLDUM
XI227 VSS WL[28] FRAM512_BITCELLDUM
XI228 VSS WL[27] FRAM512_BITCELLDUM
XI229 VSS WL[26] FRAM512_BITCELLDUM
XI230 VSS WL[25] FRAM512_BITCELLDUM
XI231 VSS WL[24] FRAM512_BITCELLDUM
XI232 VSS WL[23] FRAM512_BITCELLDUM
XI233 VSS WL[22] FRAM512_BITCELLDUM
XI234 VSS WL[21] FRAM512_BITCELLDUM
XI235 VSS WL[20] FRAM512_BITCELLDUM
XI236 VSS WL[19] FRAM512_BITCELLDUM
XI237 VSS WL[18] FRAM512_BITCELLDUM
XI238 VSS WL[17] FRAM512_BITCELLDUM
XI239 VSS WL[16] FRAM512_BITCELLDUM
XI240 VSS WL[15] FRAM512_BITCELLDUM
XI241 VSS WL[14] FRAM512_BITCELLDUM
XI242 VSS WL[13] FRAM512_BITCELLDUM
XI243 VSS WL[12] FRAM512_BITCELLDUM
XI244 VSS WL[11] FRAM512_BITCELLDUM
XI245 VSS WL[10] FRAM512_BITCELLDUM
XI246 VSS WL[9] FRAM512_BITCELLDUM
XI247 VSS WL[8] FRAM512_BITCELLDUM
XI248 VSS WL[7] FRAM512_BITCELLDUM
XI249 VSS WL[6] FRAM512_BITCELLDUM
XI250 VSS WL[5] FRAM512_BITCELLDUM
XI251 VSS WL[4] FRAM512_BITCELLDUM
XI252 VSS WL[3] FRAM512_BITCELLDUM
XI253 VSS STWL[3] FRAM512_BITCELLDUM
XI254 VSS WL[2] FRAM512_BITCELLDUM
XI255 VSS STWL[2] FRAM512_BITCELLDUM
XI256 VSS WL[1] FRAM512_BITCELLDUM
XI257 VSS STWL[1] FRAM512_BITCELLDUM
XI258 VSS WL[0] FRAM512_BITCELLDUM
XI259 VSS STWL[0] FRAM512_BITCELLDUM
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_YMX2W_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_YMX2W_FLT BLW[1] BLW[0] BLXW[1] BLXW[0] CTRCLKW CTRCLKWX DATA VDD VSS YXW[1] YXW[0]
M0 4 DATA VDD VDD P18 L=1.8E-07 W=4E-07
M1 VDD YXW[0] 3 VDD P18 L=1.8E-07 W=8E-07
M2 8 4 VDD VDD P18 L=5E-07 W=4E-07
M3 34 5 VDD VDD P18 L=1.8E-07 W=2.2E-07
M4 BLW[0] 3 VDD VDD P18 L=1.8E-07 W=1.5E-06
M5 10 CTRCLKWX 34 VDD P18 L=1.8E-07 W=2.2E-07
M6 BLXW[0] 3 BLW[0] VDD P18 L=1.8E-07 W=1.5E-06
M7 VDD 8 9 VDD P18 L=1.8E-07 W=1.2E-06
M8 VDD 3 BLXW[0] VDD P18 L=1.8E-07 W=1.5E-06
M9 25 9 VDD VDD P18 L=1.8E-07 W=1.2E-06
M10 5 10 VDD VDD P18 L=1.8E-07 W=1.6E-06
M11 BLW[0] 3 VDD VDD P18 L=1.8E-07 W=1.5E-06
M12 VDD 11 25 VDD P18 L=1.8E-07 W=1.2E-06
M13 BLXW[0] 3 BLW[0] VDD P18 L=1.8E-07 W=1.5E-06
M14 25 CTRCLKW 10 VDD P18 L=1.8E-07 W=1.2E-06
M15 VDD 3 BLXW[0] VDD P18 L=1.8E-07 W=1.5E-06
M16 26 11 VDD VDD P18 L=1.8E-07 W=1.2E-06
M17 BLXW[1] 18 VDD VDD P18 L=1.8E-07 W=1.5E-06
M18 VDD 13 26 VDD P18 L=1.8E-07 W=1.2E-06
M19 14 CTRCLKW 26 VDD P18 L=1.8E-07 W=1.2E-06
M20 BLW[1] 18 BLXW[1] VDD P18 L=1.8E-07 W=1.5E-06
M21 13 9 VDD VDD P18 L=1.8E-07 W=8E-07
M22 VDD 18 BLW[1] VDD P18 L=1.8E-07 W=1.5E-06
M23 VDD 14 12 VDD P18 L=1.8E-07 W=1.6E-06
M24 BLXW[1] 18 VDD VDD P18 L=1.8E-07 W=1.5E-06
M25 VDD VSS 16 VDD P18 L=1.8E-07 W=4E-07
M26 BLW[1] 18 BLXW[1] VDD P18 L=1.8E-07 W=1.5E-06
M27 35 CTRCLKWX 14 VDD P18 L=1.8E-07 W=2.2E-07
M28 17 16 VDD VDD P18 L=5E-07 W=4E-07
M29 VDD 18 BLW[1] VDD P18 L=1.8E-07 W=1.5E-06
M30 VDD 12 35 VDD P18 L=1.8E-07 W=2.2E-07
M31 18 YXW[1] VDD VDD P18 L=1.8E-07 W=8E-07
M32 VDD 17 11 VDD P18 L=1.8E-07 W=1.2E-06
M33 4 DATA VSS VSS N18 L=1.8E-07 W=4E-07
M34 VSS YXW[0] 3 VSS N18 L=1.8E-07 W=8E-07
M35 8 4 VSS VSS N18 L=5E-07 W=4E-07
M36 BLW[0] 5 22 VSS N18 L=1.8E-07 W=1.75E-06
M37 30 5 VSS VSS N18 L=1.8E-07 W=2.2E-07
M38 22 5 BLW[0] VSS N18 L=1.8E-07 W=1.75E-06
M39 10 CTRCLKW 30 VSS N18 L=1.8E-07 W=2.2E-07
M40 VSS 8 9 VSS N18 L=1.8E-07 W=1.2E-06
M41 VSS 3 22 VSS N18 L=1.8E-07 W=1.75E-06
M42 31 9 VSS VSS N18 L=1.8E-07 W=1.2E-06
M43 22 3 VSS VSS N18 L=1.8E-07 W=1.75E-06
M44 5 10 VSS VSS N18 L=1.8E-07 W=1.6E-06
M45 25 11 31 VSS N18 L=1.8E-07 W=1.2E-06
M46 BLXW[0] 12 22 VSS N18 L=1.8E-07 W=1.75E-06
M47 22 12 BLXW[0] VSS N18 L=1.8E-07 W=1.75E-06
M48 25 CTRCLKWX 10 VSS N18 L=1.8E-07 W=1.2E-06
M49 32 11 26 VSS N18 L=1.8E-07 W=1.2E-06
M50 VSS 13 32 VSS N18 L=1.8E-07 W=1.2E-06
M51 14 CTRCLKWX 26 VSS N18 L=1.8E-07 W=1.2E-06
M52 BLXW[1] 12 27 VSS N18 L=1.8E-07 W=1.75E-06
M53 13 9 VSS VSS N18 L=1.8E-07 W=8E-07
M54 27 12 BLXW[1] VSS N18 L=1.8E-07 W=1.75E-06
M55 VSS 14 12 VSS N18 L=1.8E-07 W=1.6E-06
M56 VSS 18 27 VSS N18 L=1.8E-07 W=1.75E-06
M57 VSS VSS 16 VSS N18 L=1.8E-07 W=4E-07
M58 27 18 VSS VSS N18 L=1.8E-07 W=1.75E-06
M59 33 CTRCLKW 14 VSS N18 L=1.8E-07 W=2.2E-07
M60 17 16 VSS VSS N18 L=5E-07 W=4E-07
M61 BLW[1] 5 27 VSS N18 L=1.8E-07 W=1.75E-06
M62 VSS 12 33 VSS N18 L=1.8E-07 W=2.2E-07
M63 27 5 BLW[1] VSS N18 L=1.8E-07 W=1.75E-06
M64 18 YXW[1] VSS VSS N18 L=1.8E-07 W=8E-07
M65 VSS 17 11 VSS N18 L=1.8E-07 W=1.2E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_YMX2R_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_YMX2R_FLT BL[1] BL[0] BLX[1] BLX[0] DOUT VDD VSS YXR[1] YXR[0] CK1 CK4
M0 BL[0] 4 23 VDD P18 L=1.8E-07 W=5E-07
M1 23 6 3 VDD P18 L=1.8E-07 W=1.4E-06
M2 VDD 3 5 VDD P18 L=2E-07 W=5.35E-07
M3 23 1 VDD VDD P18 L=1.8E-07 W=1E-06
M4 VDD 4 2 VDD P18 L=1.8E-07 W=6.7E-07
M5 23 4 BL[0] VDD P18 L=1.8E-07 W=5E-07
M6 3 6 23 VDD P18 L=1.8E-07 W=1.4E-06
M7 BL[0] 2 VDD VDD P18 L=1.8E-07 W=1E-06
M8 5 3 VDD VDD P18 L=2E-07 W=5.35E-07
M9 26 1 23 VDD P18 L=1.8E-07 W=1E-06
M10 2 4 VDD VDD P18 L=1.8E-07 W=6.7E-07
M11 BL[0] 4 23 VDD P18 L=1.8E-07 W=5E-07
M12 23 6 3 VDD P18 L=1.8E-07 W=1.4E-06
M13 BLX[0] 2 BL[0] VDD P18 L=1.8E-07 W=1E-06
M14 VDD 3 5 VDD P18 L=2E-07 W=5.35E-07
M15 VDD 1 26 VDD P18 L=1.8E-07 W=1E-06
M16 VDD 4 2 VDD P18 L=1.8E-07 W=6.7E-07
M17 VDD 2 BLX[0] VDD P18 L=1.8E-07 W=1E-06
M18 23 1 VDD VDD P18 L=1.8E-07 W=1E-06
M19 3 5 VDD VDD P18 L=2E-07 W=5.35E-07
M20 4 8 VDD VDD P18 L=1.8E-07 W=7E-07
M21 26 4 BLX[0] VDD P18 L=1.8E-07 W=5E-07
M22 5 6 26 VDD P18 L=1.8E-07 W=1.4E-06
M23 BL[0] 2 VDD VDD P18 L=1.8E-07 W=1E-06
M24 26 1 23 VDD P18 L=1.8E-07 W=1E-06
M25 VDD 5 3 VDD P18 L=2E-07 W=5.35E-07
M26 VDD 8 4 VDD P18 L=1.8E-07 W=7E-07
M27 BLX[0] 4 26 VDD P18 L=1.8E-07 W=5E-07
M28 26 6 5 VDD P18 L=1.8E-07 W=1.4E-06
M29 BLX[0] 2 BL[0] VDD P18 L=1.8E-07 W=1E-06
M30 VDD 1 26 VDD P18 L=1.8E-07 W=1E-06
M31 3 5 VDD VDD P18 L=2E-07 W=5.35E-07
M32 26 4 BLX[0] VDD P18 L=1.8E-07 W=5E-07
M33 8 YXR[0] VDD VDD P18 L=1.8E-07 W=4E-07
M34 5 6 26 VDD P18 L=1.8E-07 W=1.4E-06
M35 VDD 2 BLX[0] VDD P18 L=1.8E-07 W=1E-06
M36 13 CK4 VDD VDD P18 L=1.8E-07 W=4E-07
M37 BLX[1] 20 VDD VDD P18 L=1.8E-07 W=1E-06
M38 VDD CK1 13 VDD P18 L=1.8E-07 W=4E-07
M39 VDD YXR[1] 14 VDD P18 L=1.8E-07 W=4E-07
M40 BLX[1] 17 26 VDD P18 L=1.8E-07 W=5E-07
M41 BL[1] 20 BLX[1] VDD P18 L=1.8E-07 W=1E-06
M42 16 5 VDD VDD P18 L=1.8E-07 W=1.5E-06
M43 6 13 VDD VDD P18 L=1.8E-07 W=1.2E-06
M44 26 17 BLX[1] VDD P18 L=1.8E-07 W=5E-07
M45 17 14 VDD VDD P18 L=1.8E-07 W=7E-07
M46 VDD 20 BL[1] VDD P18 L=1.8E-07 W=1E-06
M47 VDD 15 16 VDD P18 L=1.8E-07 W=1.5E-06
M48 BLX[1] 17 26 VDD P18 L=1.8E-07 W=5E-07
M49 VDD 14 17 VDD P18 L=1.8E-07 W=7E-07
M50 BLX[1] 20 VDD VDD P18 L=1.8E-07 W=1E-06
M51 15 16 VDD VDD P18 L=1.8E-07 W=1.5E-06
M52 VDD 18 1 VDD P18 L=1.8E-07 W=1.6E-06
M53 20 17 VDD VDD P18 L=1.8E-07 W=6.7E-07
M54 BL[1] 20 BLX[1] VDD P18 L=1.8E-07 W=1E-06
M55 VDD 3 15 VDD P18 L=1.8E-07 W=1.5E-06
M56 18 CK4 VDD VDD P18 L=1.8E-07 W=4E-07
M57 23 17 BL[1] VDD P18 L=1.8E-07 W=5E-07
M58 VDD 17 20 VDD P18 L=1.8E-07 W=6.7E-07
M59 VDD 20 BL[1] VDD P18 L=1.8E-07 W=1E-06
M60 BL[1] 17 23 VDD P18 L=1.8E-07 W=5E-07
M61 VDD CK1 19 VDD P18 L=1.8E-07 W=4E-07
M62 20 17 VDD VDD P18 L=1.8E-07 W=6.7E-07
M63 DOUT 15 VDD VDD P18 L=1.8E-07 W=2E-06
M64 23 17 BL[1] VDD P18 L=1.8E-07 W=5E-07
M65 7 19 VDD VDD P18 L=1.8E-07 W=1.2E-06
M66 VDD 15 DOUT VDD P18 L=1.8E-07 W=2E-06
M67 5 3 24 VSS N18 L=2E-07 W=3E-06
M68 31 7 24 VSS N18 L=1.8E-07 W=2E-06
M69 VSS 1 31 VSS N18 L=1.8E-07 W=2E-06
M70 VSS 4 2 VSS N18 L=1.8E-07 W=6.7E-07
M71 24 3 5 VSS N18 L=2E-07 W=3E-06
M72 2 4 VSS VSS N18 L=1.8E-07 W=6.7E-07
M73 3 5 24 VSS N18 L=2E-07 W=3E-06
M74 VSS 4 2 VSS N18 L=1.8E-07 W=6.7E-07
M75 24 5 3 VSS N18 L=2E-07 W=3E-06
M76 4 8 VSS VSS N18 L=1.8E-07 W=6E-07
M77 VSS 8 4 VSS N18 L=1.8E-07 W=6E-07
M78 8 YXR[0] VSS VSS N18 L=1.8E-07 W=4E-07
M79 32 CK4 13 VSS N18 L=1.8E-07 W=4E-07
M80 VSS CK1 32 VSS N18 L=1.8E-07 W=4E-07
M81 VSS YXR[1] 14 VSS N18 L=1.8E-07 W=4E-07
M82 6 13 VSS VSS N18 L=1.8E-07 W=1.2E-06
M83 33 5 16 VSS N18 L=1.8E-07 W=1.5E-06
M84 17 14 VSS VSS N18 L=1.8E-07 W=6E-07
M85 VSS 15 33 VSS N18 L=1.8E-07 W=1.5E-06
M86 VSS 14 17 VSS N18 L=1.8E-07 W=6E-07
M87 34 16 VSS VSS N18 L=1.8E-07 W=1.5E-06
M88 VSS 18 1 VSS N18 L=1.8E-07 W=1.2E-06
M89 20 17 VSS VSS N18 L=1.8E-07 W=6.7E-07
M90 15 3 34 VSS N18 L=1.8E-07 W=1.5E-06
M91 18 CK4 VSS VSS N18 L=1.8E-07 W=8E-07
M92 VSS 17 20 VSS N18 L=1.8E-07 W=6.7E-07
M93 VSS CK1 19 VSS N18 L=1.8E-07 W=4E-07
M94 20 17 VSS VSS N18 L=1.8E-07 W=6.7E-07
M95 DOUT 15 VSS VSS N18 L=1.8E-07 W=1E-06
M96 7 19 VSS VSS N18 L=1.8E-07 W=1.2E-06
M97 VSS 15 DOUT VSS N18 L=1.8E-07 W=1E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_YMX2SAWR_AB
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_YMX2SAWR_AB BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] CK1 CK4
+CTRCLK CTRCLKX DATA QA VDD VSS YXR[1] YXR[0] YXW[1] YXW[0]
XYMUXW BLB[1] BLB[0] BLXB[1] BLXB[0] CTRCLK CTRCLKX DATA VDD VSS YXW[1] YXW[0] 
+ / FRAM512_YMX2W_FLT
XYMUXR BLA[1] BLA[0] BLXA[1] BLXA[0] QA VDD VSS YXR[1] YXR[0] CK1 CK4 / 
+ FRAM512_YMX2R_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL8T
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL8T BA BB BXA BXB VDD VSS WLA WLB
MM0 BCN BC VSS VSS N18 W=705.00N L=180.00N M=1
MM4 BB WLB BC VSS N18 W=220.00N L=225.00N M=1
MM1 BC BCN VSS VSS N18 W=705.00N L=180.00N M=1
MM2 BXA WLA BCN VSS N18 W=220.00N L=225.00N M=1
MM3 BA WLA BC VSS N18 W=220.00N L=225.00N M=1
MM7 BXB WLB BCN VSS N18 W=220.00N L=225.00N M=1
MM5 BCN BC VDD VDD P18 W=220.000N L=200.00N M=1
MM6 BC BCN VDD VDD P18 W=220.000N L=200.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL2X2
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL2X2 BA[1] BA[0] BB[1] BB[0] BXA[1] BXA[0] BXB[1] BXB[0] VDD VSS
+WLA[1] WLA[0] WLB[1] WLB[0]
XI8 BA[0] BB[0] BXA[0] BXB[0] VDD VSS WLA[0] WLB[0] FRAM512_BITCELL8T
XI11 BA[1] BB[1] BXA[1] BXB[1] VDD VSS WLA[1] WLB[1] FRAM512_BITCELL8T
XI9 BA[0] BB[0] BXA[0] BXB[0] VDD VSS WLA[1] WLB[1] FRAM512_BITCELL8T
XI10 BA[1] BB[1] BXA[1] BXB[1] VDD VSS WLA[0] WLB[0] FRAM512_BITCELL8T
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL32X2N
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL32X2N BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[31] WLA[30] WLB[31] WLB[30] FRAM512_BITCELL2X2
XI1 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[29] WLA[28] WLB[29] WLB[28] FRAM512_BITCELL2X2
XI2 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[27] WLA[26] WLB[27] WLB[26] FRAM512_BITCELL2X2
XI3 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[25] WLA[24] WLB[25] WLB[24] FRAM512_BITCELL2X2
XI4 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[23] WLA[22] WLB[23] WLB[22] FRAM512_BITCELL2X2
XI5 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[21] WLA[20] WLB[21] WLB[20] FRAM512_BITCELL2X2
XI6 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[19] WLA[18] WLB[19] WLB[18] FRAM512_BITCELL2X2
XI7 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[17] WLA[16] WLB[17] WLB[16] FRAM512_BITCELL2X2
XI8 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[15] WLA[14] WLB[15] WLB[14] FRAM512_BITCELL2X2
XI9 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[13] WLA[12] WLB[13] WLB[12] FRAM512_BITCELL2X2
XI10 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[11] WLA[10] WLB[11] WLB[10] FRAM512_BITCELL2X2
XI11 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[9] WLA[8] WLB[9] WLB[8] FRAM512_BITCELL2X2
XI12 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[7] WLA[6] WLB[7] WLB[6] FRAM512_BITCELL2X2
XI13 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[5] WLA[4] WLB[5] WLB[4] FRAM512_BITCELL2X2
XI14 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[3] WLA[2] WLB[3] WLB[2] FRAM512_BITCELL2X2
XI15 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[1] WLA[0] WLB[1] WLB[0] FRAM512_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL256X2
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL256X2 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216]
+WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206]
+WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196]
+WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126]
+WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116]
+WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106]
+WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96]
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252]
+WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242]
+WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232]
+WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222]
+WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212]
+WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202]
+WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192]
+WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182]
+WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172]
+WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162]
+WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152]
+WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142]
+WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132]
+WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122]
+WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112]
+WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102]
+WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92]
+WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82]
+WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72]
+WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] FRAM512_BITCELL32X2N
XI1 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] FRAM512_BITCELL32X2N
XI2 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] FRAM512_BITCELL32X2N
XI3 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120]
+WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110]
+WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100]
+WLB[99] WLB[98] WLB[97] WLB[96] FRAM512_BITCELL32X2N
XI4 BLXA[1] BLXA[0] BLXB[1] BLXB[0] BLA[1] BLA[0] BLB[1] BLB[0] VDD VSS
+WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150]
+WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140]
+WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130]
+WLA[129] WLA[128] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152]
+WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142]
+WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132]
+WLB[131] WLB[130] WLB[129] WLB[128] FRAM512_BITCELL32X2N
XI5 BLXA[1] BLXA[0] BLXB[1] BLXB[0] BLA[1] BLA[0] BLB[1] BLB[0] VDD VSS
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] FRAM512_BITCELL32X2N
XI6 BLXA[1] BLXA[0] BLXB[1] BLXB[0] BLA[1] BLA[0] BLB[1] BLB[0] VDD VSS
+WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214]
+WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204]
+WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194]
+WLA[193] WLA[192] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216]
+WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206]
+WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196]
+WLB[195] WLB[194] WLB[193] WLB[192] FRAM512_BITCELL32X2N
XI7 BLXA[1] BLXA[0] BLXB[1] BLXB[0] BLA[1] BLA[0] BLB[1] BLB[0] VDD VSS
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] FRAM512_BITCELL32X2N
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL2X2_STWL
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL2X2_STWL BA0 BXA0 VDD VSS WLA[3] WLA[2] WLA[1] WLA[0] WLB[3] WLB[2] WLB[1] WLB[0]
XI8 BA0 NET54 BXA0 NET53 VDD VSS WLA[0] WLB[0] FRAM512_BITCELL8T
XI11 BA3 NET46 BXA3 NET45 VDD VSS WLA[3] WLB[3] FRAM512_BITCELL8T
XI9 NET64 NET54 NET63 NET53 VDD VSS WLA[1] WLB[1] FRAM512_BITCELL8T
XI10 NET64 NET46 NET63 NET45 VDD VSS WLA[2] WLB[2] FRAM512_BITCELL8T
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL256X2ABR
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL256X2ABR BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] RDWLA[3] RDWLA[2]
+RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] VDD VSS WLA[255] WLA[254]
+WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244]
+WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234]
+WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224]
+WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214]
+WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204]
+WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194]
+WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184]
+WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174]
+WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164]
+WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154]
+WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144]
+WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134]
+WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124]
+WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114]
+WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104]
+WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94]
+WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84]
+WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74]
+WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64]
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250]
+WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240]
+WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230]
+WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220]
+WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210]
+WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200]
+WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190]
+WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180]
+WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170]
+WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160]
+WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150]
+WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140]
+WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130]
+WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120]
+WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110]
+WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100]
+WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90]
+WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80]
+WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70]
+WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216]
+WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206]
+WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196]
+WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126]
+WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116]
+WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106]
+WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96]
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252]
+WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242]
+WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232]
+WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222]
+WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212]
+WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202]
+WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192]
+WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182]
+WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172]
+WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162]
+WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152]
+WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142]
+WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132]
+WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122]
+WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112]
+WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102]
+WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92]
+WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82]
+WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72]
+WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0] FRAM512_BITCELL256X2
XI1 BLA[1] BLXA[1] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] FRAM512_BITCELL2X2_STWL
XI2 BLA[0] BLXA[0] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] FRAM512_BITCELL2X2_STWL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_ARRAY_X256Y2D1
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_ARRAY_X256Y2D1 CLKB CLKXB DATAB DOUTA RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] SACK1A SACK4A
+CLKB CLKXB DATAB DOUTA VDD VSS YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_YMX2SAWR_AB
XI1 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VSS VSS
+VSS VSS RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] VDD VSS WLA[255] WLA[254]
+WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244]
+WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234]
+WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224]
+WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214]
+WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204]
+WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194]
+WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184]
+WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174]
+WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164]
+WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154]
+WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144]
+WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134]
+WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124]
+WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114]
+WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104]
+WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94]
+WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84]
+WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74]
+WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64]
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250]
+WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240]
+WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230]
+WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220]
+WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210]
+WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200]
+WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190]
+WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180]
+WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170]
+WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160]
+WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150]
+WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140]
+WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130]
+WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120]
+WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110]
+WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100]
+WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90]
+WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80]
+WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70]
+WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] FRAM512_BITCELL256X2ABR
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_BITCELL256X2ABR_MID
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_BITCELL256X2ABR_MID BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] RDWLA[3] RDWLA[2]
+RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216]
+WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206]
+WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196]
+WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126]
+WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116]
+WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106]
+WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96]
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252]
+WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242]
+WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232]
+WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222]
+WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212]
+WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202]
+WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192]
+WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182]
+WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172]
+WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162]
+WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152]
+WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142]
+WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132]
+WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122]
+WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112]
+WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102]
+WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92]
+WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82]
+WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72]
+WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0] FRAM512_BITCELL256X2
XI1 BLA[1] BLXA[1] VDD VSS RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] FRAM512_BITCELL2X2_STWL
XI2 BLA[0] BLXA[0] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] FRAM512_BITCELL2X2_STWL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_ARRAY_X256Y2D1_MD
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_ARRAY_X256Y2D1_MD CLKB CLKXB DATAB DOUTA RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2]
+RDWLB_MID[1] RDWLB_MID[0] SACK1A SACK4A VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0]
+YXB[1] YXB[0]
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] SACK1A SACK4A
+CLKB CLKXB DATAB DOUTA VDD VSS YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_YMX2SAWR_AB
XI1 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VSS VSS
+VSS VSS VSS VSS VSS VSS RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] FRAM512_BITCELL256X2ABR_MID
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_ARRAY_X256Y2D24_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_ARRAY_X256Y2D24_RIGHT CLKB CLKXB DATAB[23] DATAB[22] DATAB[21] DATAB[20] DATAB[19] DATAB[18] DATAB[17] DATAB[16]
+DATAB[15] DATAB[14] DATAB[13] DATAB[12] DATAB[11] DATAB[10] DATAB[9] DATAB[8] DATAB[7] DATAB[6]
+DATAB[5] DATAB[4] DATAB[3] DATAB[2] DATAB[1] DATAB[0] DBL DOUTA[23] DOUTA[22] DOUTA[21]
+DOUTA[20] DOUTA[19] DOUTA[18] DOUTA[17] DOUTA[16] DOUTA[15] DOUTA[14] DOUTA[13] DOUTA[12] DOUTA[11]
+DOUTA[10] DOUTA[9] DOUTA[8] DOUTA[7] DOUTA[6] DOUTA[5] DOUTA[4] DOUTA[3] DOUTA[2] DOUTA[1]
+DOUTA[0] SACK1A SACK4A STWLA VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0]
+YXB[1] YXB[0]
XI0 DBL VDD VSS FRAM512_BITCELL_EDGE256
XI1 VSS VSS VSS VSS VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251]
+WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241]
+WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231]
+WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221]
+WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211]
+WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201]
+WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191]
+WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181]
+WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171]
+WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161]
+WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151]
+WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141]
+WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131]
+WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121]
+WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111]
+WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101]
+WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91]
+WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81]
+WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71]
+WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41]
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31]
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1]
+WLA[0] FRAM512_PCAP_DUMMY256
XI2 CLKB CLKXB DATAB[23] DOUTA[23] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI3 CLKB CLKXB DATAB[22] DOUTA[22] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI4 CLKB CLKXB DATAB[21] DOUTA[21] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI5 CLKB CLKXB DATAB[20] DOUTA[20] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI6 CLKB CLKXB DATAB[19] DOUTA[19] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI7 CLKB CLKXB DATAB[18] DOUTA[18] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI8 CLKB CLKXB DATAB[17] DOUTA[17] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI9 CLKB CLKXB DATAB[16] DOUTA[16] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI10 CLKB CLKXB DATAB[15] DOUTA[15] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI11 CLKB CLKXB DATAB[14] DOUTA[14] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI12 CLKB CLKXB DATAB[13] DOUTA[13] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI13 CLKB CLKXB DATAB[12] DOUTA[12] VSS VSS VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI14 CLKB CLKXB DATAB[11] DOUTA[11] VSS STWLA STWLA VSS VSS STWLA
+STWLA VSS SACK1A SACK4A VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0]
+YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1_MD
XI15 CLKB CLKXB DATAB[10] DOUTA[10] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI16 CLKB CLKXB DATAB[9] DOUTA[9] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI17 CLKB CLKXB DATAB[8] DOUTA[8] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI18 CLKB CLKXB DATAB[7] DOUTA[7] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI19 CLKB CLKXB DATAB[6] DOUTA[6] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI20 CLKB CLKXB DATAB[5] DOUTA[5] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI21 CLKB CLKXB DATAB[4] DOUTA[4] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI22 CLKB CLKXB DATAB[3] DOUTA[3] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI23 CLKB CLKXB DATAB[2] DOUTA[2] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI24 CLKB CLKXB DATAB[1] DOUTA[1] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI25 CLKB CLKXB DATAB[0] DOUTA[0] VSS STWLA STWLA VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_ARRAY_X256Y2D24_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_ARRAY_X256Y2D24_LEFT CLKB CLKXB DATAB[23] DATAB[22] DATAB[21] DATAB[20] DATAB[19] DATAB[18] DATAB[17] DATAB[16]
+DATAB[15] DATAB[14] DATAB[13] DATAB[12] DATAB[11] DATAB[10] DATAB[9] DATAB[8] DATAB[7] DATAB[6]
+DATAB[5] DATAB[4] DATAB[3] DATAB[2] DATAB[1] DATAB[0] DBL DOUTA[23] DOUTA[22] DOUTA[21]
+DOUTA[20] DOUTA[19] DOUTA[18] DOUTA[17] DOUTA[16] DOUTA[15] DOUTA[14] DOUTA[13] DOUTA[12] DOUTA[11]
+DOUTA[10] DOUTA[9] DOUTA[8] DOUTA[7] DOUTA[6] DOUTA[5] DOUTA[4] DOUTA[3] DOUTA[2] DOUTA[1]
+DOUTA[0] SACK1A SACK4A STWLA VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0]
+YXB[1] YXB[0]
XI0 DBL VDD VSS FRAM512_BITCELL_EDGE256
XI1 VSS VSS VSS VSS VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251]
+WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241]
+WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231]
+WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221]
+WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211]
+WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201]
+WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191]
+WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181]
+WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171]
+WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161]
+WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151]
+WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141]
+WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131]
+WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121]
+WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111]
+WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101]
+WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91]
+WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81]
+WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71]
+WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41]
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31]
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1]
+WLA[0] FRAM512_PCAP_DUMMY256
XI2 CLKB CLKXB DATAB[23] DOUTA[23] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI3 CLKB CLKXB DATAB[22] DOUTA[22] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI4 CLKB CLKXB DATAB[21] DOUTA[21] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI5 CLKB CLKXB DATAB[20] DOUTA[20] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI6 CLKB CLKXB DATAB[19] DOUTA[19] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI7 CLKB CLKXB DATAB[18] DOUTA[18] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI8 CLKB CLKXB DATAB[17] DOUTA[17] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI9 CLKB CLKXB DATAB[16] DOUTA[16] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI10 CLKB CLKXB DATAB[15] DOUTA[15] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI11 CLKB CLKXB DATAB[14] DOUTA[14] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI12 CLKB CLKXB DATAB[13] DOUTA[13] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI13 CLKB CLKXB DATAB[12] DOUTA[12] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI14 CLKB CLKXB DATAB[11] DOUTA[11] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI15 CLKB CLKXB DATAB[10] DOUTA[10] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI16 CLKB CLKXB DATAB[9] DOUTA[9] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI17 CLKB CLKXB DATAB[8] DOUTA[8] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI18 CLKB CLKXB DATAB[7] DOUTA[7] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI19 CLKB CLKXB DATAB[6] DOUTA[6] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI20 CLKB CLKXB DATAB[5] DOUTA[5] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI21 CLKB CLKXB DATAB[4] DOUTA[4] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI22 CLKB CLKXB DATAB[3] DOUTA[3] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI23 CLKB CLKXB DATAB[2] DOUTA[2] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI24 CLKB CLKXB DATAB[1] DOUTA[1] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
XI25 CLKB CLKXB DATAB[0] DOUTA[0] VSS STWLA VSS VSS SACK1A SACK4A
+VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[1] YXA[0] YXB[1] YXB[0] FRAM512_ARRAY_X256Y2D1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_SOP_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_SOP_FLT DBLA EMCLKA S[1] S[0] STWLA VDD VSS
M0 8 EMCLKA VDD VDD P18 L=1.8E-07 W=1.6E-06
M1 VDD EMCLKA 8 VDD P18 L=1.8E-07 W=1.6E-06
M2 STWLA 8 VDD VDD P18 L=1.8E-07 W=2E-06
M3 VDD 8 STWLA VDD P18 L=1.8E-07 W=2E-06
M4 STWLA 8 VDD VDD P18 L=1.8E-07 W=2E-06
M5 VDD 8 STWLA VDD P18 L=1.8E-07 W=2E-06
M6 STWLA 8 VDD VDD P18 L=1.8E-07 W=2E-06
M7 VDD S[0] 11 VDD P18 L=1.8E-07 W=1.2E-06
M8 10 S[1] VDD VDD P18 L=1.8E-07 W=1.2E-06
M9 VDD 10 3 VDD P18 L=1.8E-07 W=1.2E-06
M10 4 10 VDD VDD P18 L=1.8E-07 W=1.2E-06
M11 VDD 11 4 VDD P18 L=1.8E-07 W=1.2E-06
M12 19 11 VDD VDD P18 L=1.8E-07 W=1.2E-06
M13 5 10 19 VDD P18 L=1.8E-07 W=1.2E-06
M14 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M15 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M16 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M17 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M18 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M19 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M20 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M21 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M22 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M23 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M24 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M25 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M26 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M27 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M28 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M29 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M30 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M31 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M32 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M33 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M34 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M35 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M36 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M37 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M38 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M39 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M40 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M41 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M42 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M43 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M44 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M45 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M46 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M47 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M48 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M49 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M50 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M51 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M52 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M53 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M54 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M55 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M56 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M57 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M58 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M59 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M60 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M61 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M62 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M63 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M64 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M65 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M66 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M67 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M68 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M69 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M70 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M71 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M72 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M73 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M74 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M75 VSS 3 13 VSS N18 L=1.8E-07 W=7.05E-07
M76 13 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M77 VSS 4 15 VSS N18 L=1.8E-07 W=7.05E-07
M78 15 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M79 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M80 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M81 VSS 5 16 VSS N18 L=1.8E-07 W=7.05E-07
M82 16 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M83 VSS VDD 17 VSS N18 L=1.8E-07 W=7.05E-07
M84 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M85 13 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M86 DBLA STWLA 13 VSS N18 L=2.25E-07 W=2.2E-07
M87 15 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M88 DBLA STWLA 15 VSS N18 L=2.25E-07 W=2.2E-07
M89 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M90 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M91 16 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M92 DBLA STWLA 16 VSS N18 L=2.25E-07 W=2.2E-07
M93 17 STWLA DBLA VSS N18 L=2.25E-07 W=2.2E-07
M94 VSS S[0] 11 VSS N18 L=1.8E-07 W=1.2E-06
M95 10 S[1] VSS VSS N18 L=1.8E-07 W=1.2E-06
M96 VSS 10 3 VSS N18 L=1.8E-07 W=1.2E-06
M97 18 10 VSS VSS N18 L=1.8E-07 W=1.2E-06
M98 4 11 18 VSS N18 L=1.8E-07 W=1.2E-06
M99 5 11 VSS VSS N18 L=1.8E-07 W=1.2E-06
M100 VSS 10 5 VSS N18 L=1.8E-07 W=1.2E-06
M101 STWLA 8 VSS VSS N18 L=1.8E-07 W=1E-06
M102 VSS 8 STWLA VSS N18 L=1.8E-07 W=1E-06
M103 STWLA 8 VSS VSS N18 L=1.8E-07 W=1E-06
M104 VSS 8 STWLA VSS N18 L=1.8E-07 W=1E-06
M105 STWLA 8 VSS VSS N18 L=1.8E-07 W=1E-06
M106 8 EMCLKA VSS VSS N18 L=1.8E-07 W=8E-07
M107 VSS EMCLKA 8 VSS N18 L=1.8E-07 W=8E-07
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_SOP_W_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_SOP_W_FLT DBLB EMCLKB S[1] S[0] VDD VSS
M0 VDD S[0] 9 VDD P18 L=1.8E-07 W=1.2E-06
M1 8 S[1] VDD VDD P18 L=1.8E-07 W=1.2E-06
M2 VDD 8 3 VDD P18 L=1.8E-07 W=1.2E-06
M3 4 8 VDD VDD P18 L=1.8E-07 W=1.2E-06
M4 VDD 9 4 VDD P18 L=1.8E-07 W=1.2E-06
M5 17 9 VDD VDD P18 L=1.8E-07 W=1.2E-06
M6 5 8 17 VDD P18 L=1.8E-07 W=1.2E-06
M7 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M8 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M9 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M10 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M11 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M12 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M13 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M14 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M15 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M16 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M17 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M18 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M19 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M20 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M21 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M22 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M23 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M24 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M25 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M26 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M27 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M28 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M29 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M30 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M31 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M32 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M33 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M34 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M35 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M36 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M37 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M38 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M39 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M40 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M41 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M42 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M43 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M44 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M45 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M46 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M47 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M48 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M49 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M50 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M51 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M52 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M53 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M54 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M55 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M56 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M57 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M58 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M59 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M60 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M61 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M62 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M63 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M64 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M65 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M66 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M67 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M68 VSS 3 11 VSS N18 L=1.8E-07 W=7.05E-07
M69 11 3 VSS VSS N18 L=1.8E-07 W=7.05E-07
M70 VSS 4 13 VSS N18 L=1.8E-07 W=7.05E-07
M71 13 4 VSS VSS N18 L=1.8E-07 W=7.05E-07
M72 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M73 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M74 VSS 5 14 VSS N18 L=1.8E-07 W=7.05E-07
M75 14 5 VSS VSS N18 L=1.8E-07 W=7.05E-07
M76 VSS VDD 15 VSS N18 L=1.8E-07 W=7.05E-07
M77 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M78 11 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M79 DBLB EMCLKB 11 VSS N18 L=2.25E-07 W=2.2E-07
M80 13 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M81 DBLB EMCLKB 13 VSS N18 L=2.25E-07 W=2.2E-07
M82 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M83 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M84 14 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M85 DBLB EMCLKB 14 VSS N18 L=2.25E-07 W=2.2E-07
M86 15 EMCLKB DBLB VSS N18 L=2.25E-07 W=2.2E-07
M87 VSS S[0] 9 VSS N18 L=1.8E-07 W=1.2E-06
M88 8 S[1] VSS VSS N18 L=1.8E-07 W=1.2E-06
M89 VSS 8 3 VSS N18 L=1.8E-07 W=1.2E-06
M90 16 8 VSS VSS N18 L=1.8E-07 W=1.2E-06
M91 4 9 16 VSS N18 L=1.8E-07 W=1.2E-06
M92 5 9 VSS VSS N18 L=1.8E-07 W=1.2E-06
M93 VSS 8 5 VSS N18 L=1.8E-07 W=1.2E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_LEAFCELL_PX4_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_LEAFCELL_PX4_FLT A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] VDD VSS
M0 19 2 VDD VDD P18 L=1.8E-07 W=1E-06
M1 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M2 3 CLK 19 VDD P18 L=1.8E-07 W=8.35E-07
M3 VDD 4 19 VDD P18 L=1.8E-07 W=1E-06
M4 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M5 19 CLK 3 VDD P18 L=1.8E-07 W=8.35E-07
M6 VDD PX[0] 3 VDD P18 L=1E-06 W=2.2E-07
M7 4 A[0] VDD VDD P18 L=1.8E-07 W=4E-07
M8 19 4 VDD VDD P18 L=1.8E-07 W=1E-06
M9 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M10 3 CLK 19 VDD P18 L=1.8E-07 W=8.35E-07
M11 VDD A[0] 4 VDD P18 L=1.8E-07 W=4E-07
M12 VDD 2 19 VDD P18 L=1.8E-07 W=1E-06
M13 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M14 20 2 VDD VDD P18 L=1.8E-07 W=1E-06
M15 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M16 9 4 VDD VDD P18 L=1.8E-07 W=4E-07
M17 10 PX[1] VDD VDD P18 L=1E-06 W=2.2E-07
M18 20 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M19 VDD 9 20 VDD P18 L=1.8E-07 W=1E-06
M20 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M21 VDD 4 9 VDD P18 L=1.8E-07 W=4E-07
M22 10 CLK 20 VDD P18 L=1.8E-07 W=8.35E-07
M23 20 9 VDD VDD P18 L=1.8E-07 W=1E-06
M24 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M25 20 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M26 VDD 2 20 VDD P18 L=1.8E-07 W=1E-06
M27 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M28 21 11 VDD VDD P18 L=1.8E-07 W=1E-06
M29 PX[2] 12 VDD VDD P18 L=1.8E-07 W=2.5E-06
M30 12 CLK 21 VDD P18 L=1.8E-07 W=8.35E-07
M31 VDD 4 21 VDD P18 L=1.8E-07 W=1E-06
M32 VDD 12 PX[2] VDD P18 L=1.8E-07 W=2.5E-06
M33 21 CLK 12 VDD P18 L=1.8E-07 W=8.35E-07
M34 VDD PX[2] 12 VDD P18 L=1E-06 W=2.2E-07
M35 2 A[1] VDD VDD P18 L=1.8E-07 W=4E-07
M36 21 4 VDD VDD P18 L=1.8E-07 W=1E-06
M37 PX[2] 12 VDD VDD P18 L=1.8E-07 W=2.5E-06
M38 12 CLK 21 VDD P18 L=1.8E-07 W=8.35E-07
M39 VDD A[1] 2 VDD P18 L=1.8E-07 W=4E-07
M40 VDD 11 21 VDD P18 L=1.8E-07 W=1E-06
M41 VDD 12 PX[2] VDD P18 L=1.8E-07 W=2.5E-06
M42 22 11 VDD VDD P18 L=1.8E-07 W=1E-06
M43 PX[3] 16 VDD VDD P18 L=1.8E-07 W=2.5E-06
M44 11 2 VDD VDD P18 L=1.8E-07 W=4E-07
M45 16 PX[3] VDD VDD P18 L=1E-06 W=2.2E-07
M46 22 CLK 16 VDD P18 L=1.8E-07 W=8.35E-07
M47 VDD 9 22 VDD P18 L=1.8E-07 W=1E-06
M48 VDD 16 PX[3] VDD P18 L=1.8E-07 W=2.5E-06
M49 VDD 2 11 VDD P18 L=1.8E-07 W=4E-07
M50 16 CLK 22 VDD P18 L=1.8E-07 W=8.35E-07
M51 22 9 VDD VDD P18 L=1.8E-07 W=1E-06
M52 PX[3] 16 VDD VDD P18 L=1.8E-07 W=2.5E-06
M53 22 CLK 16 VDD P18 L=1.8E-07 W=8.35E-07
M54 VDD 11 22 VDD P18 L=1.8E-07 W=1E-06
M55 VDD 16 PX[3] VDD P18 L=1.8E-07 W=2.5E-06
M56 23 2 VSS VSS N18 L=1.8E-07 W=1E-06
M57 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M58 19 4 23 VSS N18 L=1.8E-07 W=1E-06
M59 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M60 19 CLKX 3 VSS N18 L=1.8E-07 W=1.25E-06
M61 VSS PX[0] 3 VSS N18 L=1E-06 W=2.2E-07
M62 4 A[0] VSS VSS N18 L=1.8E-07 W=4E-07
M63 24 4 19 VSS N18 L=1.8E-07 W=1E-06
M64 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M65 3 CLKX 19 VSS N18 L=1.8E-07 W=1.25E-06
M66 VSS A[0] 4 VSS N18 L=1.8E-07 W=4E-07
M67 VSS 2 24 VSS N18 L=1.8E-07 W=1E-06
M68 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M69 25 2 VSS VSS N18 L=1.8E-07 W=1E-06
M70 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M71 9 4 VSS VSS N18 L=1.8E-07 W=4E-07
M72 10 PX[1] VSS VSS N18 L=1E-06 W=2.2E-07
M73 20 CLKX 10 VSS N18 L=1.8E-07 W=1.25E-06
M74 20 9 25 VSS N18 L=1.8E-07 W=1E-06
M75 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
M76 VSS 4 9 VSS N18 L=1.8E-07 W=4E-07
M77 10 CLKX 20 VSS N18 L=1.8E-07 W=1.25E-06
M78 26 9 20 VSS N18 L=1.8E-07 W=1E-06
M79 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M80 VSS 2 26 VSS N18 L=1.8E-07 W=1E-06
M81 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
M82 27 11 VSS VSS N18 L=1.8E-07 W=1E-06
M83 PX[2] 12 VSS VSS N18 L=1.8E-07 W=1E-06
M84 21 4 27 VSS N18 L=1.8E-07 W=1E-06
M85 VSS 12 PX[2] VSS N18 L=1.8E-07 W=1E-06
M86 21 CLKX 12 VSS N18 L=1.8E-07 W=1.25E-06
M87 VSS PX[2] 12 VSS N18 L=1E-06 W=2.2E-07
M88 2 A[1] VSS VSS N18 L=1.8E-07 W=4E-07
M89 28 4 21 VSS N18 L=1.8E-07 W=1E-06
M90 PX[2] 12 VSS VSS N18 L=1.8E-07 W=1E-06
M91 12 CLKX 21 VSS N18 L=1.8E-07 W=1.25E-06
M92 VSS A[1] 2 VSS N18 L=1.8E-07 W=4E-07
M93 VSS 11 28 VSS N18 L=1.8E-07 W=1E-06
M94 VSS 12 PX[2] VSS N18 L=1.8E-07 W=1E-06
M95 29 11 VSS VSS N18 L=1.8E-07 W=1E-06
M96 PX[3] 16 VSS VSS N18 L=1.8E-07 W=1E-06
M97 11 2 VSS VSS N18 L=1.8E-07 W=4E-07
M98 16 PX[3] VSS VSS N18 L=1E-06 W=2.2E-07
M99 22 CLKX 16 VSS N18 L=1.8E-07 W=1.25E-06
M100 22 9 29 VSS N18 L=1.8E-07 W=1E-06
M101 VSS 16 PX[3] VSS N18 L=1.8E-07 W=1E-06
M102 VSS 2 11 VSS N18 L=1.8E-07 W=4E-07
M103 16 CLKX 22 VSS N18 L=1.8E-07 W=1.25E-06
M104 30 9 22 VSS N18 L=1.8E-07 W=1E-06
M105 PX[3] 16 VSS VSS N18 L=1.8E-07 W=1E-06
M106 VSS 11 30 VSS N18 L=1.8E-07 W=1E-06
M107 VSS 16 PX[3] VSS N18 L=1.8E-07 W=1E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_LEAFCELL_PX2_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_LEAFCELL_PX2_FLT A[0] CLK CLKX PX[1] PX[0] VDD VSS
M0 12 2 VDD VDD P18 L=1.8E-07 W=1E-06
M1 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M2 3 CLK 12 VDD P18 L=1.8E-07 W=8.35E-07
M3 VDD VDD 12 VDD P18 L=1.8E-07 W=1E-06
M4 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M5 12 CLK 3 VDD P18 L=1.8E-07 W=8.35E-07
M6 VDD PX[0] 3 VDD P18 L=1E-06 W=2.2E-07
M7 2 A[0] VDD VDD P18 L=1.8E-07 W=4E-07
M8 12 VDD VDD VDD P18 L=1.8E-07 W=1E-06
M9 PX[0] 3 VDD VDD P18 L=1.8E-07 W=2.5E-06
M10 3 CLK 12 VDD P18 L=1.8E-07 W=8.35E-07
M11 VDD A[0] 2 VDD P18 L=1.8E-07 W=4E-07
M12 VDD 2 12 VDD P18 L=1.8E-07 W=1E-06
M13 VDD 3 PX[0] VDD P18 L=1.8E-07 W=2.5E-06
M14 13 8 VDD VDD P18 L=1.8E-07 W=1E-06
M15 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M16 8 2 VDD VDD P18 L=1.8E-07 W=4E-07
M17 10 PX[1] VDD VDD P18 L=1E-06 W=2.2E-07
M18 13 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M19 VDD VDD 13 VDD P18 L=1.8E-07 W=1E-06
M20 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M21 VDD 2 8 VDD P18 L=1.8E-07 W=4E-07
M22 10 CLK 13 VDD P18 L=1.8E-07 W=8.35E-07
M23 13 VDD VDD VDD P18 L=1.8E-07 W=1E-06
M24 PX[1] 10 VDD VDD P18 L=1.8E-07 W=2.5E-06
M25 13 CLK 10 VDD P18 L=1.8E-07 W=8.35E-07
M26 VDD 8 13 VDD P18 L=1.8E-07 W=1E-06
M27 VDD 10 PX[1] VDD P18 L=1.8E-07 W=2.5E-06
M28 14 2 VSS VSS N18 L=1.8E-07 W=1E-06
M29 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M30 12 VDD 14 VSS N18 L=1.8E-07 W=1E-06
M31 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M32 12 CLKX 3 VSS N18 L=1.8E-07 W=1.25E-06
M33 VSS PX[0] 3 VSS N18 L=1E-06 W=2.2E-07
M34 2 A[0] VSS VSS N18 L=1.8E-07 W=4E-07
M35 15 VDD 12 VSS N18 L=1.8E-07 W=1E-06
M36 PX[0] 3 VSS VSS N18 L=1.8E-07 W=1E-06
M37 3 CLKX 12 VSS N18 L=1.8E-07 W=1.25E-06
M38 VSS A[0] 2 VSS N18 L=1.8E-07 W=4E-07
M39 VSS 2 15 VSS N18 L=1.8E-07 W=1E-06
M40 VSS 3 PX[0] VSS N18 L=1.8E-07 W=1E-06
M41 16 8 VSS VSS N18 L=1.8E-07 W=1E-06
M42 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M43 8 2 VSS VSS N18 L=1.8E-07 W=4E-07
M44 10 PX[1] VSS VSS N18 L=1E-06 W=2.2E-07
M45 13 CLKX 10 VSS N18 L=1.8E-07 W=1.25E-06
M46 13 VDD 16 VSS N18 L=1.8E-07 W=1E-06
M47 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
M48 VSS 2 8 VSS N18 L=1.8E-07 W=4E-07
M49 10 CLKX 13 VSS N18 L=1.8E-07 W=1.25E-06
M50 17 VDD 13 VSS N18 L=1.8E-07 W=1E-06
M51 PX[1] 10 VSS VSS N18 L=1.8E-07 W=1E-06
M52 VSS 8 17 VSS N18 L=1.8E-07 W=1E-06
M53 VSS 10 PX[1] VSS N18 L=1.8E-07 W=1E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_FPREDEC_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_FPREDEC_FLT A[0] A[1] A[2] CLK CLKX FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] VDD VSS WLCKX
M0 1 A[0] VDD VDD P18 L=1.8E-07 W=8E-07
M1 31 1 VDD VDD P18 L=1.8E-07 W=1E-06
M2 FCKX[2] 4 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M3 FCKX[2] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M4 4 CLK 31 VDD P18 L=1.8E-07 W=1.6E-06
M5 VDD 5 31 VDD P18 L=1.8E-07 W=1E-06
M6 WLCKX 4 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M7 VDD 6 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M8 VDD 6 4 VDD P18 L=1E-06 W=2.2E-07
M9 31 8 VDD VDD P18 L=1.8E-07 W=1E-06
M10 FCKX[2] 4 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M11 FCKX[2] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M12 VDD 4 6 VDD P18 L=1.8E-07 W=1.6E-06
M13 WLCKX 4 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M14 VDD 6 FCKX[2] VDD P18 L=1.8E-07 W=1.25E-06
M15 9 10 VDD VDD P18 L=1.8E-07 W=1.6E-06
M16 FCKX[3] 10 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M17 FCKX[3] 9 VDD VDD P18 L=1.8E-07 W=1.25E-06
M18 10 9 VDD VDD P18 L=1E-06 W=2.2E-07
M19 VDD 8 33 VDD P18 L=1.8E-07 W=1E-06
M20 WLCKX 10 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M21 VDD 9 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M22 33 5 VDD VDD P18 L=1.8E-07 W=1E-06
M23 FCKX[3] 10 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M24 FCKX[3] 9 VDD VDD P18 L=1.8E-07 W=1.25E-06
M25 33 CLK 10 VDD P18 L=1.8E-07 W=1.6E-06
M26 VDD 11 33 VDD P18 L=1.8E-07 W=1E-06
M27 WLCKX 10 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M28 VDD 9 FCKX[3] VDD P18 L=1.8E-07 W=1.25E-06
M29 35 11 VDD VDD P18 L=1.8E-07 W=1E-06
M30 FCKX[1] 12 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M31 FCKX[1] 13 VDD VDD P18 L=1.8E-07 W=1.25E-06
M32 11 1 VDD VDD P18 L=1.8E-07 W=8E-07
M33 12 CLK 35 VDD P18 L=1.8E-07 W=1.6E-06
M34 VDD 5 35 VDD P18 L=1.8E-07 W=1E-06
M35 WLCKX 12 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M36 VDD 13 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M37 VDD 13 12 VDD P18 L=1E-06 W=2.2E-07
M38 35 14 VDD VDD P18 L=1.8E-07 W=1E-06
M39 FCKX[1] 12 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M40 FCKX[1] 13 VDD VDD P18 L=1.8E-07 W=1.25E-06
M41 14 A[1] VDD VDD P18 L=1.8E-07 W=8E-07
M42 VDD 12 13 VDD P18 L=1.8E-07 W=1.6E-06
M43 WLCKX 12 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M44 VDD 13 FCKX[1] VDD P18 L=1.8E-07 W=1.25E-06
M45 15 17 VDD VDD P18 L=1.8E-07 W=1.6E-06
M46 FCKX[0] 17 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M47 FCKX[0] 15 VDD VDD P18 L=1.8E-07 W=1.25E-06
M48 17 15 VDD VDD P18 L=1E-06 W=2.2E-07
M49 VDD 14 37 VDD P18 L=1.8E-07 W=1E-06
M50 WLCKX 17 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M51 VDD 15 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M52 37 5 VDD VDD P18 L=1.8E-07 W=1E-06
M53 FCKX[0] 17 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M54 FCKX[0] 15 VDD VDD P18 L=1.8E-07 W=1.25E-06
M55 37 CLK 17 VDD P18 L=1.8E-07 W=1.6E-06
M56 VDD 1 37 VDD P18 L=1.8E-07 W=1E-06
M57 WLCKX 17 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M58 VDD 15 FCKX[0] VDD P18 L=1.8E-07 W=1.25E-06
M59 39 1 VDD VDD P18 L=1.8E-07 W=1E-06
M60 FCKX[4] 18 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M61 FCKX[4] 20 VDD VDD P18 L=1.8E-07 W=1.25E-06
M62 18 CLK 39 VDD P18 L=1.8E-07 W=1.6E-06
M63 VDD 19 39 VDD P18 L=1.8E-07 W=1E-06
M64 WLCKX 18 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M65 VDD 20 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M66 VDD 20 18 VDD P18 L=1E-06 W=2.2E-07
M67 39 14 VDD VDD P18 L=1.8E-07 W=1E-06
M68 FCKX[4] 18 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M69 FCKX[4] 20 VDD VDD P18 L=1.8E-07 W=1.25E-06
M70 VDD 18 20 VDD P18 L=1.8E-07 W=1.6E-06
M71 WLCKX 18 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M72 VDD 20 FCKX[4] VDD P18 L=1.8E-07 W=1.25E-06
M73 8 14 VDD VDD P18 L=1.8E-07 W=8E-07
M74 21 22 VDD VDD P18 L=1.8E-07 W=1.6E-06
M75 FCKX[5] 22 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M76 FCKX[5] 21 VDD VDD P18 L=1.8E-07 W=1.25E-06
M77 22 21 VDD VDD P18 L=1E-06 W=2.2E-07
M78 VDD 14 41 VDD P18 L=1.8E-07 W=1E-06
M79 WLCKX 22 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M80 VDD 21 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M81 5 A[2] VDD VDD P18 L=1.8E-07 W=8E-07
M82 41 19 VDD VDD P18 L=1.8E-07 W=1E-06
M83 FCKX[5] 22 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M84 FCKX[5] 21 VDD VDD P18 L=1.8E-07 W=1.25E-06
M85 41 CLK 22 VDD P18 L=1.8E-07 W=1.6E-06
M86 VDD 11 41 VDD P18 L=1.8E-07 W=1E-06
M87 WLCKX 22 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M88 VDD 21 FCKX[5] VDD P18 L=1.8E-07 W=1.25E-06
M89 43 11 VDD VDD P18 L=1.8E-07 W=1E-06
M90 FCKX[7] 24 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M91 FCKX[7] 25 VDD VDD P18 L=1.8E-07 W=1.25E-06
M92 24 CLK 43 VDD P18 L=1.8E-07 W=1.6E-06
M93 VDD 19 43 VDD P18 L=1.8E-07 W=1E-06
M94 WLCKX 24 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M95 VDD 25 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M96 VDD 25 24 VDD P18 L=1E-06 W=2.2E-07
M97 43 8 VDD VDD P18 L=1.8E-07 W=1E-06
M98 FCKX[7] 24 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M99 FCKX[7] 25 VDD VDD P18 L=1.8E-07 W=1.25E-06
M100 VDD 24 25 VDD P18 L=1.8E-07 W=1.6E-06
M101 WLCKX 24 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M102 VDD 25 FCKX[7] VDD P18 L=1.8E-07 W=1.25E-06
M103 26 27 VDD VDD P18 L=1.8E-07 W=1.6E-06
M104 FCKX[6] 27 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M105 FCKX[6] 26 VDD VDD P18 L=1.8E-07 W=1.25E-06
M106 27 26 VDD VDD P18 L=1E-06 W=2.2E-07
M107 VDD 8 45 VDD P18 L=1.8E-07 W=1E-06
M108 WLCKX 27 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M109 VDD 26 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M110 45 19 VDD VDD P18 L=1.8E-07 W=1E-06
M111 FCKX[6] 27 WLCKX VDD P18 L=1.8E-07 W=1.25E-06
M112 FCKX[6] 26 VDD VDD P18 L=1.8E-07 W=1.25E-06
M113 45 CLK 27 VDD P18 L=1.8E-07 W=1.6E-06
M114 19 5 VDD VDD P18 L=1.8E-07 W=8E-07
M115 VDD 1 45 VDD P18 L=1.8E-07 W=1E-06
M116 WLCKX 27 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M117 VDD 26 FCKX[6] VDD P18 L=1.8E-07 W=1.25E-06
M118 47 1 VSS VSS N18 L=1.8E-07 W=1E-06
M119 FCKX[2] 6 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M120 4 CLKX 31 VSS N18 L=1.8E-07 W=1.6E-06
M121 48 5 47 VSS N18 L=1.8E-07 W=1E-06
M122 WLCKX 6 FCKX[2] VSS N18 L=1.8E-07 W=1.25E-06
M123 VSS 6 4 VSS N18 L=1E-06 W=2.2E-07
M124 31 8 48 VSS N18 L=1.8E-07 W=1E-06
M125 FCKX[2] 6 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M126 1 A[0] VSS VSS N18 L=1.8E-07 W=8E-07
M127 VSS 4 6 VSS N18 L=1.8E-07 W=1.6E-06
M128 WLCKX 6 FCKX[2] VSS N18 L=1.8E-07 W=1.25E-06
M129 9 10 VSS VSS N18 L=1.8E-07 W=1.6E-06
M130 FCKX[3] 9 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M131 10 9 VSS VSS N18 L=1E-06 W=2.2E-07
M132 49 8 33 VSS N18 L=1.8E-07 W=1E-06
M133 WLCKX 9 FCKX[3] VSS N18 L=1.8E-07 W=1.25E-06
M134 11 1 VSS VSS N18 L=1.8E-07 W=8E-07
M135 50 5 49 VSS N18 L=1.8E-07 W=1E-06
M136 FCKX[3] 9 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M137 33 CLKX 10 VSS N18 L=1.8E-07 W=1.6E-06
M138 VSS 11 50 VSS N18 L=1.8E-07 W=1E-06
M139 WLCKX 9 FCKX[3] VSS N18 L=1.8E-07 W=1.25E-06
M140 51 11 VSS VSS N18 L=1.8E-07 W=1E-06
M141 FCKX[1] 13 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M142 12 CLKX 35 VSS N18 L=1.8E-07 W=1.6E-06
M143 52 5 51 VSS N18 L=1.8E-07 W=1E-06
M144 WLCKX 13 FCKX[1] VSS N18 L=1.8E-07 W=1.25E-06
M145 VSS 13 12 VSS N18 L=1E-06 W=2.2E-07
M146 35 14 52 VSS N18 L=1.8E-07 W=1E-06
M147 FCKX[1] 13 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M148 VSS 12 13 VSS N18 L=1.8E-07 W=1.6E-06
M149 WLCKX 13 FCKX[1] VSS N18 L=1.8E-07 W=1.25E-06
M150 15 17 VSS VSS N18 L=1.8E-07 W=1.6E-06
M151 FCKX[0] 15 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M152 17 15 VSS VSS N18 L=1E-06 W=2.2E-07
M153 53 14 37 VSS N18 L=1.8E-07 W=1E-06
M154 WLCKX 15 FCKX[0] VSS N18 L=1.8E-07 W=1.25E-06
M155 14 A[1] VSS VSS N18 L=1.8E-07 W=8E-07
M156 54 5 53 VSS N18 L=1.8E-07 W=1E-06
M157 FCKX[0] 15 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M158 37 CLKX 17 VSS N18 L=1.8E-07 W=1.6E-06
M159 VSS 1 54 VSS N18 L=1.8E-07 W=1E-06
M160 WLCKX 15 FCKX[0] VSS N18 L=1.8E-07 W=1.25E-06
M161 55 1 VSS VSS N18 L=1.8E-07 W=1E-06
M162 FCKX[4] 20 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M163 18 CLKX 39 VSS N18 L=1.8E-07 W=1.6E-06
M164 8 14 VSS VSS N18 L=1.8E-07 W=8E-07
M165 56 19 55 VSS N18 L=1.8E-07 W=1E-06
M166 WLCKX 20 FCKX[4] VSS N18 L=1.8E-07 W=1.25E-06
M167 VSS 20 18 VSS N18 L=1E-06 W=2.2E-07
M168 39 14 56 VSS N18 L=1.8E-07 W=1E-06
M169 FCKX[4] 20 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M170 VSS 18 20 VSS N18 L=1.8E-07 W=1.6E-06
M171 WLCKX 20 FCKX[4] VSS N18 L=1.8E-07 W=1.25E-06
M172 21 22 VSS VSS N18 L=1.8E-07 W=1.6E-06
M173 FCKX[5] 21 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M174 22 21 VSS VSS N18 L=1E-06 W=2.2E-07
M175 57 14 41 VSS N18 L=1.8E-07 W=1E-06
M176 WLCKX 21 FCKX[5] VSS N18 L=1.8E-07 W=1.25E-06
M177 58 19 57 VSS N18 L=1.8E-07 W=1E-06
M178 FCKX[5] 21 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M179 41 CLKX 22 VSS N18 L=1.8E-07 W=1.6E-06
M180 VSS 11 58 VSS N18 L=1.8E-07 W=1E-06
M181 WLCKX 21 FCKX[5] VSS N18 L=1.8E-07 W=1.25E-06
M182 59 11 VSS VSS N18 L=1.8E-07 W=1E-06
M183 FCKX[7] 25 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M184 5 A[2] VSS VSS N18 L=1.8E-07 W=8E-07
M185 24 CLKX 43 VSS N18 L=1.8E-07 W=1.6E-06
M186 60 19 59 VSS N18 L=1.8E-07 W=1E-06
M187 WLCKX 25 FCKX[7] VSS N18 L=1.8E-07 W=1.25E-06
M188 VSS 25 24 VSS N18 L=1E-06 W=2.2E-07
M189 43 8 60 VSS N18 L=1.8E-07 W=1E-06
M190 FCKX[7] 25 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M191 VSS 24 25 VSS N18 L=1.8E-07 W=1.6E-06
M192 WLCKX 25 FCKX[7] VSS N18 L=1.8E-07 W=1.25E-06
M193 19 5 VSS VSS N18 L=1.8E-07 W=8E-07
M194 26 27 VSS VSS N18 L=1.8E-07 W=1.6E-06
M195 FCKX[6] 26 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M196 27 26 VSS VSS N18 L=1E-06 W=2.2E-07
M197 61 8 45 VSS N18 L=1.8E-07 W=1E-06
M198 WLCKX 26 FCKX[6] VSS N18 L=1.8E-07 W=1.25E-06
M199 62 19 61 VSS N18 L=1.8E-07 W=1E-06
M200 FCKX[6] 26 WLCKX VSS N18 L=1.8E-07 W=1.25E-06
M201 45 CLKX 27 VSS N18 L=1.8E-07 W=1.6E-06
M202 VSS 1 62 VSS N18 L=1.8E-07 W=1E-06
M203 WLCKX 26 FCKX[6] VSS N18 L=1.8E-07 W=1.25E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_YPREDEC2_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_YPREDEC2_FLT A[0] CLK CLKX VDD VSS YCKX YX[1] YX[0]
M0 13 VDD VDD VDD P18 L=1.8E-07 W=1E-06
M1 YX[0] 4 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M2 YX[0] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M3 4 CLK 13 VDD P18 L=1.8E-07 W=1.6E-06
M4 VDD 5 13 VDD P18 L=1.8E-07 W=1E-06
M5 YCKX 4 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M6 VDD 6 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M7 VDD 6 4 VDD P18 L=1E-06 W=2.2E-07
M8 YX[0] 4 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M9 YX[0] 6 VDD VDD P18 L=1.8E-07 W=1.25E-06
M10 VDD A[0] 5 VDD P18 L=1.8E-07 W=8E-07
M11 VDD 4 6 VDD P18 L=1.8E-07 W=1.6E-06
M12 YCKX 4 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M13 VDD 6 YX[0] VDD P18 L=1.8E-07 W=1.25E-06
M14 10 5 VDD VDD P18 L=1.8E-07 W=8E-07
M15 8 9 VDD VDD P18 L=1.8E-07 W=1.6E-06
M16 YX[1] 9 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M17 YX[1] 8 VDD VDD P18 L=1.8E-07 W=1.25E-06
M18 9 8 VDD VDD P18 L=1E-06 W=2.2E-07
M19 YCKX 9 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M20 VDD 8 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M21 16 10 VDD VDD P18 L=1.8E-07 W=1E-06
M22 YX[1] 9 YCKX VDD P18 L=1.8E-07 W=1.25E-06
M23 YX[1] 8 VDD VDD P18 L=1.8E-07 W=1.25E-06
M24 16 CLK 9 VDD P18 L=1.8E-07 W=1.6E-06
M25 VDD VDD 16 VDD P18 L=1.8E-07 W=1E-06
M26 YCKX 9 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M27 VDD 8 YX[1] VDD P18 L=1.8E-07 W=1.25E-06
M28 17 VDD VSS VSS N18 L=1.8E-07 W=1E-06
M29 YX[0] 6 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M30 4 CLKX 13 VSS N18 L=1.8E-07 W=1.6E-06
M31 13 5 17 VSS N18 L=1.8E-07 W=1E-06
M32 YCKX 6 YX[0] VSS N18 L=1.8E-07 W=1.25E-06
M33 VSS 6 4 VSS N18 L=1E-06 W=2.2E-07
M34 YX[0] 6 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M35 VSS A[0] 5 VSS N18 L=1.8E-07 W=8E-07
M36 VSS 4 6 VSS N18 L=1.8E-07 W=1.6E-06
M37 YCKX 6 YX[0] VSS N18 L=1.8E-07 W=1.25E-06
M38 10 5 VSS VSS N18 L=1.8E-07 W=8E-07
M39 8 9 VSS VSS N18 L=1.8E-07 W=1.6E-06
M40 YX[1] 8 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M41 9 8 VSS VSS N18 L=1E-06 W=2.2E-07
M42 YCKX 8 YX[1] VSS N18 L=1.8E-07 W=1.25E-06
M43 18 10 16 VSS N18 L=1.8E-07 W=1E-06
M44 YX[1] 8 YCKX VSS N18 L=1.8E-07 W=1.25E-06
M45 16 CLKX 9 VSS N18 L=1.8E-07 W=1.6E-06
M46 VSS VDD 18 VSS N18 L=1.8E-07 W=1E-06
M47 YCKX 8 YX[1] VSS N18 L=1.8E-07 W=1.25E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_TP_CLKW_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_TP_CLKW_FLT CEN CLK DCTRCLK DCTRCLKX EMCLKB FB INTCLKX S[0] VDD VMINE VSS
M0 6 10 VDD VDD P18 L=1.8E-07 W=4E-06
M1 VDD 10 6 VDD P18 L=1.8E-07 W=4E-06
M2 3 6 VDD VDD P18 L=1.8E-07 W=2E-06
M3 VDD 6 3 VDD P18 L=1.8E-07 W=2E-06
M4 8 2 3 VDD P18 L=1.8E-07 W=2E-06
M5 3 2 8 VDD P18 L=1.8E-07 W=2E-06
M6 VDD S[0] 7 VDD P18 L=1.8E-07 W=8E-07
M7 1 7 VDD VDD P18 L=1.8E-07 W=1.2E-06
M8 2 1 VDD VDD P18 L=1.8E-07 W=1.2E-06
M9 8 1 29 VDD P18 L=1.8E-07 W=2E-06
M10 29 1 8 VDD P18 L=1.8E-07 W=2E-06
M11 29 6 VDD VDD P18 L=1.8E-07 W=2E-06
M12 VDD 5 29 VDD P18 L=1.8E-07 W=2E-06
M13 VDD 3 5 VDD P18 L=1.8E-07 W=2E-06
M14 EMCLKB 8 VDD VDD P18 L=1.8E-07 W=4E-06
M15 VDD 8 EMCLKB VDD P18 L=1.8E-07 W=4E-06
M16 11 FB VDD VDD P18 L=1.8E-07 W=1.2E-06
M17 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M18 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M19 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M20 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M21 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M22 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M23 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M24 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M25 10 9 VDD VDD P18 L=1.8E-07 W=1E-06
M26 VDD 9 10 VDD P18 L=1.8E-07 W=1E-06
M27 VDD 15 9 VDD P18 L=1.8E-07 W=2.1E-06
M28 9 15 VDD VDD P18 L=1.8E-07 W=2.1E-06
M29 VDD 11 9 VDD P18 L=1.8E-07 W=2.1E-06
M30 9 11 VDD VDD P18 L=1.8E-07 W=2.1E-06
M31 VDD 15 35 VDD P18 L=1.8E-07 W=2E-06
M32 35 15 VDD VDD P18 L=1.8E-07 W=2E-06
M33 VDD 15 35 VDD P18 L=1.8E-07 W=2E-06
M34 35 15 VDD VDD P18 L=1.8E-07 W=2E-06
M35 VDD 15 35 VDD P18 L=1.8E-07 W=2E-06
M36 35 15 VDD VDD P18 L=1.8E-07 W=2E-06
M37 10 CLK 35 VDD P18 L=1.8E-07 W=2E-06
M38 35 CLK 10 VDD P18 L=1.8E-07 W=2E-06
M39 10 CLK 35 VDD P18 L=1.8E-07 W=2E-06
M40 35 CLK 10 VDD P18 L=1.8E-07 W=2E-06
M41 10 CLK 35 VDD P18 L=1.8E-07 W=2E-06
M42 35 CLK 10 VDD P18 L=1.8E-07 W=2E-06
M43 FB 6 VDD VDD P18 L=1.8E-07 W=2.4E-06
M44 VDD 6 FB VDD P18 L=1.8E-07 W=2.4E-06
M45 FB 6 VDD VDD P18 L=1.8E-07 W=2.4E-06
M46 17 10 VDD VDD P18 L=1.8E-07 W=9.95E-07
M47 VDD 10 17 VDD P18 L=1.8E-07 W=3.28E-06
M48 17 10 VDD VDD P18 L=1.8E-07 W=3.28E-06
M49 VDD 10 17 VDD P18 L=1.8E-07 W=3.28E-06
M50 17 10 VDD VDD P18 L=1.8E-07 W=3.28E-06
M51 15 VMINE VDD VDD P18 L=1.8E-07 W=2.8E-06
M52 42 CLK VDD VDD P18 L=1.8E-07 W=2E-06
M53 18 CEN 42 VDD P18 L=1.8E-07 W=2E-06
M54 43 16 VDD VDD P18 L=1.8E-07 W=2E-06
M55 19 CLK 43 VDD P18 L=1.8E-07 W=2E-06
M56 20 19 VDD VDD P18 L=1.8E-07 W=2E-06
M57 12 20 VDD VDD P18 L=1.8E-07 W=2E-06
M58 VDD 20 12 VDD P18 L=1.8E-07 W=2E-06
M59 12 20 VDD VDD P18 L=1.8E-07 W=2E-06
M60 VDD 16 18 VDD P18 L=1E-06 W=2.2E-07
M61 10 17 VDD VDD P18 L=1E-06 W=2.2E-07
M62 VDD CLK 21 VDD P18 L=1.8E-07 W=1.2E-06
M63 16 18 VDD VDD P18 L=1.8E-07 W=1.2E-06
M64 DCTRCLK 24 VDD VDD P18 L=1.8E-07 W=3.06E-06
M65 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=3.06E-06
M66 DCTRCLK 24 VDD VDD P18 L=1.8E-07 W=3.06E-06
M67 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=3.06E-06
M68 DCTRCLK 24 VDD VDD P18 L=1.8E-07 W=3.06E-06
M69 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=3.06E-06
M70 27 24 VDD VDD P18 L=1.8E-07 W=3E-06
M71 VDD 24 27 VDD P18 L=1.8E-07 W=3E-06
M72 24 17 38 VDD P18 L=1.8E-07 W=3.5E-06
M73 38 17 24 VDD P18 L=1.8E-07 W=3.5E-06
M74 VDD 26 38 VDD P18 L=1.8E-07 W=3.5E-06
M75 38 26 VDD VDD P18 L=1.8E-07 W=3.5E-06
M76 VDD 17 25 VDD P18 L=1.8E-07 W=5E-07
M77 VDD 24 DCTRCLK VDD P18 L=1.8E-07 W=1.66E-06
M78 VDD 17 INTCLKX VDD P18 L=1.8E-07 W=2.8E-06
M79 INTCLKX 17 VDD VDD P18 L=1.8E-07 W=2.8E-06
M80 VDD 17 INTCLKX VDD P18 L=1.8E-07 W=2.8E-06
M81 INTCLKX 17 VDD VDD P18 L=1.8E-07 W=2.8E-06
M82 VDD 17 INTCLKX VDD P18 L=1.8E-07 W=2.8E-06
M83 VDD 25 26 VDD P18 L=1.8E-07 W=5E-07
M84 DCTRCLKX 27 VDD VDD P18 L=1.8E-07 W=6.67E-06
M85 VDD 27 DCTRCLKX VDD P18 L=1.8E-07 W=6.67E-06
M86 DCTRCLKX 27 VDD VDD P18 L=1.8E-07 W=6.67E-06
M87 6 10 VSS VSS N18 L=1.8E-07 W=2E-06
M88 VSS 10 6 VSS N18 L=1.8E-07 W=2E-06
M89 3 6 VSS VSS N18 L=1.8E-07 W=2E-06
M90 VSS 6 3 VSS N18 L=1.8E-07 W=2E-06
M91 8 1 3 VSS N18 L=1.8E-07 W=2E-06
M92 3 1 8 VSS N18 L=1.8E-07 W=2E-06
M93 8 2 29 VSS N18 L=1.8E-07 W=2E-06
M94 29 2 8 VSS N18 L=1.8E-07 W=2E-06
M95 40 6 29 VSS N18 L=1.8E-07 W=2E-06
M96 VSS 5 40 VSS N18 L=1.8E-07 W=2E-06
M97 EMCLKB 8 VSS VSS N18 L=1.8E-07 W=2E-06
M98 VSS 8 EMCLKB VSS N18 L=1.8E-07 W=2E-06
M99 1 7 VSS VSS N18 L=1.8E-07 W=1.2E-06
M100 2 1 VSS VSS N18 L=1.8E-07 W=1.2E-06
M101 VSS 3 5 VSS N18 L=1.8E-07 W=1E-06
M102 VSS S[0] 7 VSS N18 L=1.8E-07 W=8E-07
M103 9 15 33 VSS N18 L=1.8E-07 W=2.1E-06
M104 33 15 9 VSS N18 L=1.8E-07 W=2.1E-06
M105 VSS 11 33 VSS N18 L=1.8E-07 W=2.1E-06
M106 33 11 VSS VSS N18 L=1.8E-07 W=2.1E-06
M107 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M108 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M109 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M110 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M111 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M112 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M113 10 CLK 34 VSS N18 L=1.8E-07 W=2.5E-06
M114 34 CLK 10 VSS N18 L=1.8E-07 W=2.5E-06
M115 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M116 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M117 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M118 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M119 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M120 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M121 VSS 12 34 VSS N18 L=1.8E-07 W=2.5E-06
M122 34 12 VSS VSS N18 L=1.8E-07 W=2.5E-06
M123 11 FB VSS VSS N18 L=1.8E-07 W=1.2E-06
M124 VSS CLK 21 VSS N18 L=1.8E-07 W=1.2E-06
M125 41 21 VSS VSS N18 L=1.8E-07 W=2E-06
M126 18 CEN 41 VSS N18 L=1.8E-07 W=2E-06
M127 16 18 VSS VSS N18 L=1.8E-07 W=1.2E-06
M128 19 16 VSS VSS N18 L=1.8E-07 W=1E-06
M129 VSS CLK 19 VSS N18 L=1.8E-07 W=1E-06
M130 20 19 VSS VSS N18 L=1.8E-07 W=1E-06
M131 12 20 VSS VSS N18 L=1.8E-07 W=1.5E-06
M132 VSS 20 12 VSS N18 L=1.8E-07 W=1.5E-06
M133 VSS 10 17 VSS N18 L=1.8E-07 W=1.75E-06
M134 17 10 VSS VSS N18 L=1.8E-07 W=1.75E-06
M135 VSS 10 17 VSS N18 L=1.8E-07 W=1.75E-06
M136 17 10 VSS VSS N18 L=1.8E-07 W=1.75E-06
M137 10 17 VSS VSS N18 L=1E-06 W=2.2E-07
M138 18 16 VSS VSS N18 L=1E-06 W=2.2E-07
M139 15 VMINE VSS VSS N18 L=1.8E-07 W=1.4E-06
M140 24 17 VSS VSS N18 L=1.8E-07 W=3.5E-06
M141 VSS 17 24 VSS N18 L=1.8E-07 W=3.5E-06
M142 24 26 VSS VSS N18 L=1.8E-07 W=3.5E-06
M143 VSS 26 24 VSS N18 L=1.8E-07 W=3.5E-06
M144 VSS 24 DCTRCLK VSS N18 L=1.8E-07 W=3.335E-06
M145 DCTRCLK 24 VSS VSS N18 L=1.8E-07 W=3.335E-06
M146 VSS 24 DCTRCLK VSS N18 L=1.8E-07 W=3.335E-06
M147 27 24 VSS VSS N18 L=1.8E-07 W=3E-06
M148 VSS 24 27 VSS N18 L=1.8E-07 W=3E-06
M149 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=4.4E-06
M150 INTCLKX 17 VSS VSS N18 L=1.8E-07 W=4.4E-06
M151 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=4.4E-06
M152 INTCLKX 17 VSS VSS N18 L=1.8E-07 W=4.4E-06
M153 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=4.4E-06
M154 INTCLKX 17 VSS VSS N18 L=1.8E-07 W=3E-06
M155 VSS 17 INTCLKX VSS N18 L=1.8E-07 W=3E-06
M156 VSS 25 26 VSS N18 L=1.8E-07 W=5E-07
M157 VSS 17 25 VSS N18 L=1.8E-07 W=5E-07
M158 DCTRCLKX 27 VSS VSS N18 L=1.8E-07 W=5E-06
M159 VSS 27 DCTRCLKX VSS N18 L=1.8E-07 W=5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_LOGIC_Y2_W_X256
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_LOGIC_Y2_W_X256 AB[8] AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CENB
+CLKB DCTRCLK DCTRCLKX EMCLKB FB FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3]
+FCKXB[2] FCKXB[1] FCKXB[0] PXAB[3] PXAB[2] PXAB[1] PXAB[0] PXBB[3] PXBB[2] PXBB[1]
+PXBB[0] PXCB[1] PXCB[0] S[0] VDD VMINE VSS YXW[1] YXW[0]
XPXB4B AB[6] AB[7] DCTRCLK DCTRCLKX PXBB[3] PXBB[2] PXBB[1] PXBB[0] VDD VSS 
+ FRAM512_LEAFCELL_PX4_FLT
XPA AB[4] AB[5] DCTRCLK DCTRCLKX PXAB[3] PXAB[2] PXAB[1] PXAB[0] VDD VSS 
+ FRAM512_LEAFCELL_PX4_FLT
XPXC2B AB[8] DCTRCLK DCTRCLKX PXCB[1] PXCB[0] VDD VSS FRAM512_LEAFCELL_PX2_FLT
XFPRE AB[1] AB[2] AB[3] DCTRCLK DCTRCLKX FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] 
+ FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0] VDD VSS INTCLKXB FRAM512_FPREDEC_FLT
XI0 AB[0] DCTRCLK DCTRCLKX VDD VSS INTCLKXB YXW[1] YXW[0] FRAM512_YPREDEC2_FLT
XCLKDRV CENB CLKB DCTRCLK DCTRCLKX EMCLKB FB INTCLKXB S[0] VDD VMINE VSS 
+ FRAM512_TP_CLKW_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_CLK_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_CLK_FLT ACTRCLK ACTRCLKX CEN CLK EMCLKA FB INTCLKX S[0] SACK1 SACK4
+VDD VMINE VSS
M0 4 VMINE VDD VDD P18 L=1.8E-07 W=2.8E-06
M1 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M2 7 2 VDD VDD P18 L=1.8E-07 W=4E-06
M3 ACTRCLKX ACTRCLK VDD VDD P18 L=1.8E-07 W=3.5E-06
M4 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M5 VDD 4 36 VDD P18 L=1.8E-07 W=2E-06
M6 VDD 2 7 VDD P18 L=1.8E-07 W=4E-06
M7 VDD ACTRCLK ACTRCLKX VDD P18 L=1.8E-07 W=3.5E-06
M8 VDD CLK 6 VDD P18 L=1.8E-07 W=1.2E-06
M9 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M10 36 4 VDD VDD P18 L=1.8E-07 W=2E-06
M11 ACTRCLKX ACTRCLK VDD VDD P18 L=1.8E-07 W=3.5E-06
M12 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M13 VDD 4 36 VDD P18 L=1.8E-07 W=2E-06
M14 47 CLK VDD VDD P18 L=1.8E-07 W=2E-06
M15 26 7 VDD VDD P18 L=1.8E-07 W=2E-06
M16 VDD ACTRCLK ACTRCLKX VDD P18 L=1.8E-07 W=3.5E-06
M17 10 CEN 47 VDD P18 L=1.8E-07 W=2E-06
M18 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M19 36 4 VDD VDD P18 L=1.8E-07 W=2E-06
M20 VDD 7 26 VDD P18 L=1.8E-07 W=2E-06
M21 ACTRCLK 11 VDD VDD P18 L=1.8E-07 W=3.5E-06
M22 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M23 VDD 4 36 VDD P18 L=1.8E-07 W=2E-06
M24 VDD 11 ACTRCLK VDD P18 L=1.8E-07 W=3.5E-06
M25 12 10 VDD VDD P18 L=1.8E-07 W=1.2E-06
M26 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M27 36 4 VDD VDD P18 L=1.8E-07 W=2E-06
M28 29 14 26 VDD P18 L=1.8E-07 W=2E-06
M29 ACTRCLK 11 VDD VDD P18 L=1.8E-07 W=3.5E-06
M30 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M31 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M32 2 CLK 36 VDD P18 L=1.8E-07 W=2E-06
M33 26 14 29 VDD P18 L=1.8E-07 W=2E-06
M34 VDD 11 ACTRCLK VDD P18 L=1.8E-07 W=3.5E-06
M35 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M36 VDD 9 INTCLKX VDD P18 L=1.8E-07 W=1.4E-06
M37 36 CLK 2 VDD P18 L=1.8E-07 W=2E-06
M38 VDD 12 10 VDD P18 L=1E-06 W=2.2E-07
M39 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M40 INTCLKX 9 VDD VDD P18 L=1.8E-07 W=1.4E-06
M41 2 CLK 36 VDD P18 L=1.8E-07 W=2E-06
M42 VDD S[0] 16 VDD P18 L=1.8E-07 W=8E-07
M43 11 9 38 VDD P18 L=1.8E-07 W=2.5E-06
M44 48 12 VDD VDD P18 L=1.8E-07 W=2E-06
M45 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M46 36 CLK 2 VDD P18 L=1.8E-07 W=2E-06
M47 38 9 11 VDD P18 L=1.8E-07 W=2.5E-06
M48 13 16 VDD VDD P18 L=1.8E-07 W=1.2E-06
M49 19 CLK 48 VDD P18 L=1.8E-07 W=2E-06
M50 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M51 2 CLK 36 VDD P18 L=1.8E-07 W=2E-06
M52 VDD 18 38 VDD P18 L=1.8E-07 W=2.5E-06
M53 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M54 36 CLK 2 VDD P18 L=1.8E-07 W=2E-06
M55 38 18 VDD VDD P18 L=1.8E-07 W=2.5E-06
M56 14 13 VDD VDD P18 L=1.8E-07 W=1.2E-06
M57 21 19 VDD VDD P18 L=1.8E-07 W=2E-06
M58 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M59 SACK1 9 VDD VDD P18 L=1.8E-07 W=1.86E-06
M60 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M61 29 13 39 VDD P18 L=1.8E-07 W=2E-06
M62 FB 7 VDD VDD P18 L=1.8E-07 W=2.4E-06
M63 VDD 9 SACK1 VDD P18 L=1.8E-07 W=3.035E-06
M64 20 21 VDD VDD P18 L=1.8E-07 W=2E-06
M65 2 17 VDD VDD P18 L=1.8E-07 W=1E-06
M66 VDD 22 18 VDD P18 L=1.8E-07 W=5E-07
M67 VDD 9 22 VDD P18 L=1.8E-07 W=5E-07
M68 39 13 29 VDD P18 L=1.8E-07 W=2E-06
M69 VDD 7 FB VDD P18 L=1.8E-07 W=2.4E-06
M70 SACK1 9 VDD VDD P18 L=1.8E-07 W=3.035E-06
M71 VDD 21 20 VDD P18 L=1.8E-07 W=2E-06
M72 VDD 17 2 VDD P18 L=1.8E-07 W=1E-06
M73 FB 7 VDD VDD P18 L=1.8E-07 W=2.4E-06
M74 VDD 9 SACK1 VDD P18 L=1.8E-07 W=3.035E-06
M75 20 21 VDD VDD P18 L=1.8E-07 W=2E-06
M76 39 7 VDD VDD P18 L=1.8E-07 W=2E-06
M77 SACK1 9 VDD VDD P18 L=1.8E-07 W=3.035E-06
M78 24 9 VDD VDD P18 L=1.8E-07 W=5E-07
M79 28 24 VDD VDD P18 L=1.8E-07 W=5E-07
M80 30 FB VDD VDD P18 L=1.8E-07 W=1.2E-06
M81 2 9 VDD VDD P18 L=1E-06 W=2.2E-07
M82 VDD 25 39 VDD P18 L=1.8E-07 W=2E-06
M83 9 2 VDD VDD P18 L=1.8E-07 W=9.95E-07
M84 VDD 27 SACK4 VDD P18 L=1.8E-07 W=2.8E-06
M85 VDD 26 25 VDD P18 L=1.8E-07 W=2E-06
M86 VDD 4 17 VDD P18 L=1.8E-07 W=2.1E-06
M87 VDD 2 9 VDD P18 L=1.8E-07 W=3.28E-06
M88 43 9 27 VDD P18 L=1.8E-07 W=3E-06
M89 SACK4 27 VDD VDD P18 L=1.8E-07 W=2.8E-06
M90 17 4 VDD VDD P18 L=1.8E-07 W=2.1E-06
M91 9 2 VDD VDD P18 L=1.8E-07 W=3.28E-06
M92 VDD 28 43 VDD P18 L=1.8E-07 W=3E-06
M93 VDD 27 SACK4 VDD P18 L=1.8E-07 W=2.8E-06
M94 EMCLKA 29 VDD VDD P18 L=1.8E-07 W=4E-06
M95 VDD 30 17 VDD P18 L=1.8E-07 W=2.1E-06
M96 VDD 2 9 VDD P18 L=1.8E-07 W=3.28E-06
M97 43 28 VDD VDD P18 L=1.8E-07 W=3E-06
M98 SACK4 27 VDD VDD P18 L=1.8E-07 W=2.8E-06
M99 VDD 29 EMCLKA VDD P18 L=1.8E-07 W=4E-06
M100 17 30 VDD VDD P18 L=1.8E-07 W=2.1E-06
M101 9 2 VDD VDD P18 L=1.8E-07 W=3.28E-06
M102 27 9 43 VDD P18 L=1.8E-07 W=3E-06
M103 VDD 27 SACK4 VDD P18 L=1.8E-07 W=2.8E-06
M104 4 VMINE VSS VSS N18 L=1.8E-07 W=1.4E-06
M105 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M106 7 2 VSS VSS N18 L=1.8E-07 W=2E-06
M107 ACTRCLKX ACTRCLK VSS VSS N18 L=1.8E-07 W=1.75E-06
M108 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M109 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M110 VSS 2 7 VSS N18 L=1.8E-07 W=2E-06
M111 VSS ACTRCLK ACTRCLKX VSS N18 L=1.8E-07 W=1.75E-06
M112 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M113 VSS CLK 6 VSS N18 L=1.8E-07 W=1.2E-06
M114 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M115 ACTRCLKX ACTRCLK VSS VSS N18 L=1.8E-07 W=1.75E-06
M116 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M117 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M118 45 6 VSS VSS N18 L=1.8E-07 W=2E-06
M119 26 7 VSS VSS N18 L=1.8E-07 W=2E-06
M120 VSS ACTRCLK ACTRCLKX VSS N18 L=1.8E-07 W=1.75E-06
M121 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M122 10 CEN 45 VSS N18 L=1.8E-07 W=2E-06
M123 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M124 VSS 7 26 VSS N18 L=1.8E-07 W=2E-06
M125 ACTRCLK 11 VSS VSS N18 L=1.8E-07 W=1.75E-06
M126 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M127 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M128 VSS 11 ACTRCLK VSS N18 L=1.8E-07 W=1.75E-06
M129 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M130 12 10 VSS VSS N18 L=1.8E-07 W=1.2E-06
M131 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M132 29 13 26 VSS N18 L=1.8E-07 W=2E-06
M133 ACTRCLK 11 VSS VSS N18 L=1.8E-07 W=1.75E-06
M134 2 CLK 35 VSS N18 L=1.8E-07 W=2.5E-06
M135 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M136 26 13 29 VSS N18 L=1.8E-07 W=2E-06
M137 VSS 11 ACTRCLK VSS N18 L=1.8E-07 W=1.75E-06
M138 35 CLK 2 VSS N18 L=1.8E-07 W=2.5E-06
M139 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M140 10 12 VSS VSS N18 L=1E-06 W=2.2E-07
M141 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M142 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M143 VSS S[0] 16 VSS N18 L=1.8E-07 W=8E-07
M144 11 9 VSS VSS N18 L=1.8E-07 W=2.5E-06
M145 19 12 VSS VSS N18 L=1.8E-07 W=1E-06
M146 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M147 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=2.1E-06
M148 VSS 9 11 VSS N18 L=1.8E-07 W=2.5E-06
M149 13 16 VSS VSS N18 L=1.8E-07 W=1.2E-06
M150 VSS CLK 19 VSS N18 L=1.8E-07 W=1E-06
M151 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M152 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=2.1E-06
M153 11 18 VSS VSS N18 L=1.8E-07 W=2.5E-06
M154 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M155 VSS 9 INTCLKX VSS N18 L=1.8E-07 W=1.4E-06
M156 VSS 18 11 VSS N18 L=1.8E-07 W=2.5E-06
M157 14 13 VSS VSS N18 L=1.8E-07 W=1.2E-06
M158 21 19 VSS VSS N18 L=1.8E-07 W=1E-06
M159 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M160 INTCLKX 9 VSS VSS N18 L=1.8E-07 W=1.4E-06
M161 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M162 29 14 39 VSS N18 L=1.8E-07 W=2E-06
M163 20 21 VSS VSS N18 L=1.8E-07 W=1.5E-06
M164 VSS 20 35 VSS N18 L=1.8E-07 W=2.5E-06
M165 VSS 22 18 VSS N18 L=1.8E-07 W=5E-07
M166 VSS 9 22 VSS N18 L=1.8E-07 W=5E-07
M167 39 14 29 VSS N18 L=1.8E-07 W=2E-06
M168 SACK1 9 VSS VSS N18 L=1.8E-07 W=1.75E-06
M169 VSS 21 20 VSS N18 L=1.8E-07 W=1.5E-06
M170 35 20 VSS VSS N18 L=1.8E-07 W=2.5E-06
M171 VSS 9 SACK1 VSS N18 L=1.8E-07 W=1.75E-06
M172 2 9 VSS VSS N18 L=1E-06 W=2.2E-07
M173 46 7 39 VSS N18 L=1.8E-07 W=2E-06
M174 SACK1 9 VSS VSS N18 L=1.8E-07 W=1.75E-06
M175 24 9 VSS VSS N18 L=1.8E-07 W=5E-07
M176 28 24 VSS VSS N18 L=1.8E-07 W=5E-07
M177 30 FB VSS VSS N18 L=1.8E-07 W=1.2E-06
M178 VSS 25 46 VSS N18 L=1.8E-07 W=2E-06
M179 VSS 9 SACK1 VSS N18 L=1.8E-07 W=1.75E-06
M180 VSS 26 25 VSS N18 L=1.8E-07 W=1E-06
M181 17 4 42 VSS N18 L=1.8E-07 W=2.1E-06
M182 VSS 2 9 VSS N18 L=1.8E-07 W=1.75E-06
M183 27 9 VSS VSS N18 L=1.8E-07 W=1.5E-06
M184 SACK4 27 VSS VSS N18 L=1.8E-07 W=1.75E-06
M185 42 4 17 VSS N18 L=1.8E-07 W=2.1E-06
M186 9 2 VSS VSS N18 L=1.8E-07 W=1.75E-06
M187 VSS 28 27 VSS N18 L=1.8E-07 W=1.5E-06
M188 VSS 27 SACK4 VSS N18 L=1.8E-07 W=1.75E-06
M189 EMCLKA 29 VSS VSS N18 L=1.8E-07 W=2E-06
M190 VSS 30 42 VSS N18 L=1.8E-07 W=2.1E-06
M191 VSS 2 9 VSS N18 L=1.8E-07 W=1.75E-06
M192 27 28 VSS VSS N18 L=1.8E-07 W=1.5E-06
M193 SACK4 27 VSS VSS N18 L=1.8E-07 W=1.75E-06
M194 VSS 29 EMCLKA VSS N18 L=1.8E-07 W=2E-06
M195 42 30 VSS VSS N18 L=1.8E-07 W=2.1E-06
M196 9 2 VSS VSS N18 L=1.8E-07 W=1.75E-06
M197 VSS 9 27 VSS N18 L=1.8E-07 W=1.5E-06
M198 VSS 27 SACK4 VSS N18 L=1.8E-07 W=1.75E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_LOGIC_Y2_R_X256
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_LOGIC_Y2_R_X256 AA[8] AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] CENA
+CLKA EMCLKA FB FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1]
+FCKXA[0] PXAA[3] PXAA[2] PXAA[1] PXAA[0] PXBA[3] PXBA[2] PXBA[1] PXBA[0] PXCA[1]
+PXCA[0] S[0] SACK1 SACK4 VDD VMINE VSS YXR[1] YXR[0]
XPXB4A AA[6] AA[7] ACTRCLK ACTRCLKX PXBA[3] PXBA[2] PXBA[1] PXBA[0] VDD VSS 
+ FRAM512_LEAFCELL_PX4_FLT
XPA AA[4] AA[5] ACTRCLK ACTRCLKX PXAA[3] PXAA[2] PXAA[1] PXAA[0] VDD VSS 
+ FRAM512_LEAFCELL_PX4_FLT
XPXC2A AA[8] ACTRCLK ACTRCLKX PXCA[1] PXCA[0] VDD VSS FRAM512_LEAFCELL_PX2_FLT
XFPRE AA[1] AA[2] AA[3] ACTRCLK ACTRCLKX FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] 
+ FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0] VDD VSS INTCLKXA FRAM512_FPREDEC_FLT
XI0 AA[0] ACTRCLK ACTRCLKX VDD VSS INTCLKXA YXR[1] YXR[0] FRAM512_YPREDEC2_FLT
XCLKDRV ACTRCLK ACTRCLKX CENA CLKA EMCLKA FB INTCLKXA S[0] SACK1 SACK4 VDD 
+ VMINE VSS FRAM512_CLK_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_XDEC_FLT
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_XDEC_FLT FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA PXB
+PXC VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
M0 6 4 VDD VDD P18 L=1.8E-07 W=1E-06
M1 VDD 4 6 VDD P18 L=1.8E-07 W=1E-06
M2 4 5 VDD VDD P18 L=1.8E-07 W=1.5E-06
M3 VDD 5 4 VDD P18 L=1.8E-07 W=1.5E-06
M4 VDD PXA 5 VDD P18 L=1.8E-07 W=1E-06
M5 5 PXB VDD VDD P18 L=1.8E-07 W=1E-06
M6 VDD PXC 5 VDD P18 L=1.8E-07 W=1E-06
M7 VDD 4 7 VDD P18 L=1.8E-07 W=1E-06
M8 8 4 VDD VDD P18 L=1.8E-07 W=1E-06
M9 VDD 4 9 VDD P18 L=1.8E-07 W=1E-06
M10 10 4 VDD VDD P18 L=1.8E-07 W=1E-06
M11 VDD 4 11 VDD P18 L=1.8E-07 W=1E-06
M12 12 4 VDD VDD P18 L=1.8E-07 W=1E-06
M13 VDD 4 13 VDD P18 L=1.8E-07 W=1E-06
M14 14 4 VDD VDD P18 L=1.8E-07 W=1E-06
M15 7 6 FCKX[0] VDD P18 L=1.8E-07 W=8E-07
M16 FCKX[1] 6 8 VDD P18 L=1.8E-07 W=8E-07
M17 9 6 FCKX[2] VDD P18 L=1.8E-07 W=8E-07
M18 FCKX[3] 6 10 VDD P18 L=1.8E-07 W=8E-07
M19 11 6 FCKX[4] VDD P18 L=1.8E-07 W=8E-07
M20 FCKX[5] 6 12 VDD P18 L=1.8E-07 W=8E-07
M21 13 6 FCKX[6] VDD P18 L=1.8E-07 W=8E-07
M22 FCKX[7] 6 14 VDD P18 L=1.8E-07 W=8E-07
M23 15 7 VDD VDD P18 L=1.8E-07 W=8E-07
M24 VDD 7 15 VDD P18 L=1.8E-07 W=8E-07
M25 16 8 VDD VDD P18 L=1.8E-07 W=8E-07
M26 VDD 8 16 VDD P18 L=1.8E-07 W=8E-07
M27 17 9 VDD VDD P18 L=1.8E-07 W=8E-07
M28 VDD 9 17 VDD P18 L=1.8E-07 W=8E-07
M29 18 10 VDD VDD P18 L=1.8E-07 W=8E-07
M30 VDD 10 18 VDD P18 L=1.8E-07 W=8E-07
M31 19 11 VDD VDD P18 L=1.8E-07 W=8E-07
M32 VDD 11 19 VDD P18 L=1.8E-07 W=8E-07
M33 20 12 VDD VDD P18 L=1.8E-07 W=8E-07
M34 VDD 12 20 VDD P18 L=1.8E-07 W=8E-07
M35 21 13 VDD VDD P18 L=1.8E-07 W=8E-07
M36 VDD 13 21 VDD P18 L=1.8E-07 W=8E-07
M37 22 14 VDD VDD P18 L=1.8E-07 W=8E-07
M38 VDD 14 22 VDD P18 L=1.8E-07 W=8E-07
M39 23 15 VDD VDD P18 L=1.8E-07 W=2E-06
M40 VDD 15 23 VDD P18 L=1.8E-07 W=2E-06
M41 24 16 VDD VDD P18 L=1.8E-07 W=2E-06
M42 VDD 16 24 VDD P18 L=1.8E-07 W=2E-06
M43 25 17 VDD VDD P18 L=1.8E-07 W=2E-06
M44 VDD 17 25 VDD P18 L=1.8E-07 W=2E-06
M45 26 18 VDD VDD P18 L=1.8E-07 W=2E-06
M46 VDD 18 26 VDD P18 L=1.8E-07 W=2E-06
M47 27 19 VDD VDD P18 L=1.8E-07 W=2E-06
M48 VDD 19 27 VDD P18 L=1.8E-07 W=2E-06
M49 28 20 VDD VDD P18 L=1.8E-07 W=2E-06
M50 VDD 20 28 VDD P18 L=1.8E-07 W=2E-06
M51 29 21 VDD VDD P18 L=1.8E-07 W=2E-06
M52 VDD 21 29 VDD P18 L=1.8E-07 W=2E-06
M53 30 22 VDD VDD P18 L=1.8E-07 W=2E-06
M54 VDD 22 30 VDD P18 L=1.8E-07 W=2E-06
M55 WL[0] 23 VDD VDD P18 L=1.8E-07 W=7E-06
M56 VDD 23 WL[0] VDD P18 L=1.8E-07 W=7E-06
M57 WL[1] 24 VDD VDD P18 L=1.8E-07 W=7E-06
M58 VDD 24 WL[1] VDD P18 L=1.8E-07 W=7E-06
M59 WL[2] 25 VDD VDD P18 L=1.8E-07 W=7E-06
M60 VDD 25 WL[2] VDD P18 L=1.8E-07 W=7E-06
M61 WL[3] 26 VDD VDD P18 L=1.8E-07 W=7E-06
M62 VDD 26 WL[3] VDD P18 L=1.8E-07 W=7E-06
M63 WL[4] 27 VDD VDD P18 L=1.8E-07 W=7E-06
M64 VDD 27 WL[4] VDD P18 L=1.8E-07 W=7E-06
M65 WL[5] 28 VDD VDD P18 L=1.8E-07 W=7E-06
M66 VDD 28 WL[5] VDD P18 L=1.8E-07 W=7E-06
M67 WL[6] 29 VDD VDD P18 L=1.8E-07 W=7E-06
M68 VDD 29 WL[6] VDD P18 L=1.8E-07 W=7E-06
M69 WL[7] 30 VDD VDD P18 L=1.8E-07 W=7E-06
M70 VDD 30 WL[7] VDD P18 L=1.8E-07 W=7E-06
M71 78 PXA 5 VSS N18 L=1.8E-07 W=1.6E-06
M72 79 PXB 78 VSS N18 L=1.8E-07 W=1.6E-06
M73 VSS PXC 79 VSS N18 L=1.8E-07 W=1.6E-06
M74 6 4 VSS VSS N18 L=1.8E-07 W=1E-06
M75 VSS 4 6 VSS N18 L=1.8E-07 W=1E-06
M76 4 5 VSS VSS N18 L=1.8E-07 W=1E-06
M77 VSS 5 4 VSS N18 L=1.8E-07 W=1E-06
M78 7 4 FCKX[0] VSS N18 L=1.8E-07 W=1E-06
M79 FCKX[1] 4 8 VSS N18 L=1.8E-07 W=1E-06
M80 9 4 FCKX[2] VSS N18 L=1.8E-07 W=1E-06
M81 FCKX[3] 4 10 VSS N18 L=1.8E-07 W=1E-06
M82 11 4 FCKX[4] VSS N18 L=1.8E-07 W=1E-06
M83 FCKX[5] 4 12 VSS N18 L=1.8E-07 W=1E-06
M84 13 4 FCKX[6] VSS N18 L=1.8E-07 W=1E-06
M85 FCKX[7] 4 14 VSS N18 L=1.8E-07 W=1E-06
M86 15 7 VSS VSS N18 L=1.8E-07 W=4E-07
M87 VSS 7 15 VSS N18 L=1.8E-07 W=4E-07
M88 16 8 VSS VSS N18 L=1.8E-07 W=4E-07
M89 VSS 8 16 VSS N18 L=1.8E-07 W=4E-07
M90 17 9 VSS VSS N18 L=1.8E-07 W=4E-07
M91 VSS 9 17 VSS N18 L=1.8E-07 W=4E-07
M92 18 10 VSS VSS N18 L=1.8E-07 W=4E-07
M93 VSS 10 18 VSS N18 L=1.8E-07 W=4E-07
M94 19 11 VSS VSS N18 L=1.8E-07 W=4E-07
M95 VSS 11 19 VSS N18 L=1.8E-07 W=4E-07
M96 20 12 VSS VSS N18 L=1.8E-07 W=4E-07
M97 VSS 12 20 VSS N18 L=1.8E-07 W=4E-07
M98 21 13 VSS VSS N18 L=1.8E-07 W=4E-07
M99 VSS 13 21 VSS N18 L=1.8E-07 W=4E-07
M100 22 14 VSS VSS N18 L=1.8E-07 W=4E-07
M101 VSS 14 22 VSS N18 L=1.8E-07 W=4E-07
M102 23 15 VSS VSS N18 L=1.8E-07 W=1.2E-06
M103 VSS 15 23 VSS N18 L=1.8E-07 W=1.2E-06
M104 24 16 VSS VSS N18 L=1.8E-07 W=1.2E-06
M105 VSS 16 24 VSS N18 L=1.8E-07 W=1.2E-06
M106 25 17 VSS VSS N18 L=1.8E-07 W=1.2E-06
M107 VSS 17 25 VSS N18 L=1.8E-07 W=1.2E-06
M108 26 18 VSS VSS N18 L=1.8E-07 W=1.2E-06
M109 VSS 18 26 VSS N18 L=1.8E-07 W=1.2E-06
M110 27 19 VSS VSS N18 L=1.8E-07 W=1.2E-06
M111 VSS 19 27 VSS N18 L=1.8E-07 W=1.2E-06
M112 28 20 VSS VSS N18 L=1.8E-07 W=1.2E-06
M113 VSS 20 28 VSS N18 L=1.8E-07 W=1.2E-06
M114 29 21 VSS VSS N18 L=1.8E-07 W=1.2E-06
M115 VSS 21 29 VSS N18 L=1.8E-07 W=1.2E-06
M116 30 22 VSS VSS N18 L=1.8E-07 W=1.2E-06
M117 VSS 22 30 VSS N18 L=1.8E-07 W=1.2E-06
M118 WL[0] 23 VSS VSS N18 L=1.8E-07 W=3.5E-06
M119 VSS 23 WL[0] VSS N18 L=1.8E-07 W=3.5E-06
M120 WL[1] 24 VSS VSS N18 L=1.8E-07 W=3.5E-06
M121 VSS 24 WL[1] VSS N18 L=1.8E-07 W=3.5E-06
M122 WL[2] 25 VSS VSS N18 L=1.8E-07 W=3.5E-06
M123 VSS 25 WL[2] VSS N18 L=1.8E-07 W=3.5E-06
M124 WL[3] 26 VSS VSS N18 L=1.8E-07 W=3.5E-06
M125 VSS 26 WL[3] VSS N18 L=1.8E-07 W=3.5E-06
M126 WL[4] 27 VSS VSS N18 L=1.8E-07 W=3.5E-06
M127 VSS 27 WL[4] VSS N18 L=1.8E-07 W=3.5E-06
M128 WL[5] 28 VSS VSS N18 L=1.8E-07 W=3.5E-06
M129 VSS 28 WL[5] VSS N18 L=1.8E-07 W=3.5E-06
M130 WL[6] 29 VSS VSS N18 L=1.8E-07 W=3.5E-06
M131 VSS 29 WL[6] VSS N18 L=1.8E-07 W=3.5E-06
M132 WL[7] 30 VSS VSS N18 L=1.8E-07 W=3.5E-06
M133 VSS 30 WL[7] VSS N18 L=1.8E-07 W=3.5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512_XDEC32
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512_XDEC32 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2]
+PXA[1] PXA[0] PXB[3] PXB[2] PXB[1] PXB[0] PXC[1] PXC[0] VDD VSS
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[3]
+PXC[1] VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249]
+WL[248] FRAM512_XDEC_FLT
XI1 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[3]
+PXC[1] VDD VSS WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] FRAM512_XDEC_FLT
XI2 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[1] VDD VSS WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] FRAM512_XDEC_FLT
XI3 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[1] VDD VSS WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] FRAM512_XDEC_FLT
XI4 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[2]
+PXC[1] VDD VSS WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217]
+WL[216] FRAM512_XDEC_FLT
XI5 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[2]
+PXC[1] VDD VSS WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209]
+WL[208] FRAM512_XDEC_FLT
XI6 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[1] VDD VSS WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] FRAM512_XDEC_FLT
XI7 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[1] VDD VSS WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] FRAM512_XDEC_FLT
XI8 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[1] VDD VSS WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] FRAM512_XDEC_FLT
XI9 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[1] VDD VSS WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177]
+WL[176] FRAM512_XDEC_FLT
XI10 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[1] VDD VSS WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169]
+WL[168] FRAM512_XDEC_FLT
XI11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[1] VDD VSS WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] FRAM512_XDEC_FLT
XI12 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[1] VDD VSS WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] FRAM512_XDEC_FLT
XI13 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[1] VDD VSS WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] FRAM512_XDEC_FLT
XI14 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[1] VDD VSS WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137]
+WL[136] FRAM512_XDEC_FLT
XI15 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[1] VDD VSS WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129]
+WL[128] FRAM512_XDEC_FLT
XI16 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[3]
+PXC[0] VDD VSS WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] FRAM512_XDEC_FLT
XI17 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[3]
+PXC[0] VDD VSS WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] FRAM512_XDEC_FLT
XI18 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[0] VDD VSS WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] FRAM512_XDEC_FLT
XI19 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[0] VDD VSS WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97]
+WL[96] FRAM512_XDEC_FLT
XI20 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[2]
+PXC[0] VDD VSS WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89]
+WL[88] FRAM512_XDEC_FLT
XI21 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[2]
+PXC[0] VDD VSS WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] FRAM512_XDEC_FLT
XI22 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[0] VDD VSS WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] FRAM512_XDEC_FLT
XI23 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[0] VDD VSS WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] FRAM512_XDEC_FLT
XI24 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[0] VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] FRAM512_XDEC_FLT
XI25 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[0] VDD VSS WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] FRAM512_XDEC_FLT
XI26 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[0] VDD VSS WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] FRAM512_XDEC_FLT
XI27 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[0] VDD VSS WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] FRAM512_XDEC_FLT
XI28 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[0] VDD VSS WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] FRAM512_XDEC_FLT
XI29 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[0] VDD VSS WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] FRAM512_XDEC_FLT
XI30 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[0] VDD VSS WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] FRAM512_XDEC_FLT
XI31 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[0] VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0] FRAM512_XDEC_FLT
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    FRAM512
* View Name:    schematic
************************************************************************

.SUBCKT FRAM512 AA[8] AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] AB[8]
+AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CENA CENB
+CLKA CLKB DB[47] DB[46] DB[45] DB[44] DB[43] DB[42] DB[41] DB[40]
+DB[39] DB[38] DB[37] DB[36] DB[35] DB[34] DB[33] DB[32] DB[31] DB[30]
+DB[29] DB[28] DB[27] DB[26] DB[25] DB[24] DB[23] DB[22] DB[21] DB[20]
+DB[19] DB[18] DB[17] DB[16] DB[15] DB[14] DB[13] DB[12] DB[11] DB[10]
+DB[9] DB[8] DB[7] DB[6] DB[5] DB[4] DB[3] DB[2] DB[1] DB[0]
+QA[47] QA[46] QA[45] QA[44] QA[43] QA[42] QA[41] QA[40] QA[39] QA[38]
+QA[37] QA[36] QA[35] QA[34] QA[33] QA[32] QA[31] QA[30] QA[29] QA[28]
+QA[27] QA[26] QA[25] QA[24] QA[23] QA[22] QA[21] QA[20] QA[19] QA[18]
+QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] QA[11] QA[10] QA[9] QA[8]
+QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] VDD VSS
XI0 DCTRCLK DCTRCLKX DB[47] DB[46] DB[45] DB[44] DB[43] DB[42] DB[41] DB[40]
+DB[39] DB[38] DB[37] DB[36] DB[35] DB[34] DB[33] DB[32] DB[31] DB[30]
+DB[29] DB[28] DB[27] DB[26] DB[25] DB[24] DBLA QA[47] QA[46] QA[45]
+QA[44] QA[43] QA[42] QA[41] QA[40] QA[39] QA[38] QA[37] QA[36] QA[35]
+QA[34] QA[33] QA[32] QA[31] QA[30] QA[29] QA[28] QA[27] QA[26] QA[25]
+QA[24] SACK1 SACK4 STWLA VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] YXR[1] YXR[0]
+YXW[1] YXW[0] FRAM512_ARRAY_X256Y2D24_RIGHT
XI1 DCTRCLK DCTRCLKX DB[23] DB[22] DB[21] DB[20] DB[19] DB[18] DB[17] DB[16]
+DB[15] DB[14] DB[13] DB[12] DB[11] DB[10] DB[9] DB[8] DB[7] DB[6]
+DB[5] DB[4] DB[3] DB[2] DB[1] DB[0] DBLB QA[23] QA[22] QA[21]
+QA[20] QA[19] QA[18] QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] QA[11]
+QA[10] QA[9] QA[8] QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1]
+QA[0] SACK1 SACK4 STWLA VDD VSS WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] YXR[1] YXR[0]
+YXW[1] YXW[0] FRAM512_ARRAY_X256Y2D24_LEFT
XI2 DBLA EMCLKA VSS VDD STWLA VDD VSS FRAM512_SOP_FLT
XI3 DBLB EMCLKB VSS VDD VDD VSS FRAM512_SOP_W_FLT
XI4 AB[8] AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CENB
+CLKB DCTRCLK DCTRCLKX EMCLKB DBLB FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3]
+FCKXB[2] FCKXB[1] FCKXB[0] PXAB[3] PXAB[2] PXAB[1] PXAB[0] PXBB[3] PXBB[2] PXBB[1]
+PXBB[0] PXCB[1] PXCB[0] VSS VDD VSS VSS YXW[1] YXW[0] FRAM512_LOGIC_Y2_W_X256
XI5 AA[8] AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] CENA
+CLKA EMCLKA DBLA FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1]
+FCKXA[0] PXAA[3] PXAA[2] PXAA[1] PXAA[0] PXBA[3] PXBA[2] PXBA[1] PXBA[0] PXCA[1]
+PXCA[0] VSS SACK1 SACK4 VDD VSS VSS YXR[1] YXR[0] FRAM512_LOGIC_Y2_R_X256
XI6 FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0] PXAB[3] PXAB[2]
+PXAB[1] PXAB[0] PXBB[3] PXBB[2] PXBB[1] PXBB[0] PXCB[1] PXCB[0] VDD VSS
+WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246]
+WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236]
+WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226]
+WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216]
+WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206]
+WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196]
+WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186]
+WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176]
+WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166]
+WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156]
+WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146]
+WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136]
+WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126]
+WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116]
+WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106]
+WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96]
+WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86]
+WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76]
+WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66]
+WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] FRAM512_XDEC32
XI7 FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0] PXAA[3] PXAA[2]
+PXAA[1] PXAA[0] PXBA[3] PXBA[2] PXBA[1] PXBA[0] PXCA[1] PXCA[0] VDD VSS
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216]
+WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206]
+WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196]
+WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126]
+WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116]
+WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106]
+WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96]
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] FRAM512_XDEC32
.ENDS
