#     Copyright (c) 2022 SMIC                                                       
#     Filename:      RAM512.lef                                                   
#     IP code:       S018RF2P                                                         
#     Version:       0.2.b                                                        
#     CreateDate:    Mon Oct 31 21:43:20 CST 2022                                                     
                    
#    LEF for 2-PORT Register File                                                               
#    SMIC 0.18um G Logic Process                                                       
#    Configuration: -instname RAM512 -rows 128 -bits 24 -mux 4  



# DISCLAIMER                                                                           #
#                                                                                      #  
#   SMIC hereby provides the quality information to you but makes no claims,           #
# promises or guarantees about the accuracy, completeness, or adequacy of the          #
# information herein. The information contained herein is provided on an "AS IS"       #
# basis without any warranty, and SMIC assumes no obligation to provide support        #
# of any kind or otherwise maintain the information.                                   #  
#   SMIC disclaims any representation that the information does not infringe any       #
# intellectual property rights or proprietary rights of any third parties. SMIC        #
# makes no other warranty, whether express, implied or statutory as to any             #
# matter whatsoever, including but not limited to the accuracy or sufficiency of       #
# any information or the merchantability and fitness for a particular purpose.         #
# Neither SMIC nor any of its representatives shall be liable for any cause of         #
# action incurred to connect to this service.                                          #  
#                                                                                      #
# STATEMENT OF USE AND CONFIDENTIALITY                                                 #  
#                                                                                      #  
#   The following/attached material contains confidential and proprietary              #  
# information of SMIC. This material is based upon information which SMIC              #  
# considers reliable, but SMIC neither represents nor warrants that such               #
# information is accurate or complete, and it must not be relied upon as such.         #
# This information was prepared for informational purposes and is for the use          #
# by SMIC's customer only. SMIC reserves the right to make changes in the              #  
# information at any time without notice.                                              #  
#   No part of this information may be reproduced, transmitted, transcribed,           #  
# stored in a retrieval system, or translated into any human or computer               # 
# language, in any form or by any means, electronic, mechanical, magnetic,             #  
# optical, chemical, manual, or otherwise, without the prior written consent of        #
# SMIC. Any unauthorized use or disclosure of this material is strictly                #  
# prohibited and may be unlawful. By accepting this material, the receiving            #  
# party shall be deemed to have acknowledged, accepted, and agreed to be bound         #
# by the foregoing limitations and restrictions. Thank you.                            #  
#                                                                                      #  


MACRO RAM512
CLASS BLOCK ;
ORIGIN 0 0 ;
SIZE 676.66 BY 272.265 ;
SYMMETRY X Y R90 ;

PIN QA[11]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 8.905 271.625 9.975 272.265 ;
LAYER METAL2 ;
RECT 8.905 271.625 9.975 272.265 ;
LAYER METAL3 ;
RECT 8.905 271.625 9.975 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[11]

PIN DB[11]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL2 ;
RECT 18.725 0.0 19.795 0.64 ;
LAYER METAL3 ;
RECT 18.725 0.0 19.795 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[11]

PIN QA[10]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 32.145 271.625 33.215 272.265 ;
LAYER METAL2 ;
RECT 32.145 271.625 33.215 272.265 ;
LAYER METAL3 ;
RECT 32.145 271.625 33.215 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[10]

PIN DB[10]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL2 ;
RECT 41.965 0.0 43.035 0.64 ;
LAYER METAL3 ;
RECT 41.965 0.0 43.035 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[10]

PIN QA[9]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 55.385 271.625 56.455 272.265 ;
LAYER METAL2 ;
RECT 55.385 271.625 56.455 272.265 ;
LAYER METAL3 ;
RECT 55.385 271.625 56.455 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[9]

PIN DB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL2 ;
RECT 65.205 0.0 66.275 0.64 ;
LAYER METAL3 ;
RECT 65.205 0.0 66.275 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[9]

PIN QA[8]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 78.625 271.625 79.695 272.265 ;
LAYER METAL2 ;
RECT 78.625 271.625 79.695 272.265 ;
LAYER METAL3 ;
RECT 78.625 271.625 79.695 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[8]

PIN DB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL2 ;
RECT 88.445 0.0 89.515 0.64 ;
LAYER METAL3 ;
RECT 88.445 0.0 89.515 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[8]

PIN QA[7]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 101.865 271.625 102.935 272.265 ;
LAYER METAL2 ;
RECT 101.865 271.625 102.935 272.265 ;
LAYER METAL3 ;
RECT 101.865 271.625 102.935 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[7]

PIN DB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL2 ;
RECT 111.685 0.0 112.755 0.64 ;
LAYER METAL3 ;
RECT 111.685 0.0 112.755 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[7]

PIN QA[6]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 125.105 271.625 126.175 272.265 ;
LAYER METAL2 ;
RECT 125.105 271.625 126.175 272.265 ;
LAYER METAL3 ;
RECT 125.105 271.625 126.175 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[6]

PIN DB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL2 ;
RECT 134.925 0.0 135.995 0.64 ;
LAYER METAL3 ;
RECT 134.925 0.0 135.995 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[6]

PIN QA[5]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 148.345 271.625 149.415 272.265 ;
LAYER METAL2 ;
RECT 148.345 271.625 149.415 272.265 ;
LAYER METAL3 ;
RECT 148.345 271.625 149.415 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[5]

PIN DB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL2 ;
RECT 158.165 0.0 159.235 0.64 ;
LAYER METAL3 ;
RECT 158.165 0.0 159.235 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[5]

PIN QA[4]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 171.585 271.625 172.655 272.265 ;
LAYER METAL2 ;
RECT 171.585 271.625 172.655 272.265 ;
LAYER METAL3 ;
RECT 171.585 271.625 172.655 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[4]

PIN DB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL2 ;
RECT 181.405 0.0 182.475 0.64 ;
LAYER METAL3 ;
RECT 181.405 0.0 182.475 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[4]

PIN QA[3]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 194.825 271.625 195.895 272.265 ;
LAYER METAL2 ;
RECT 194.825 271.625 195.895 272.265 ;
LAYER METAL3 ;
RECT 194.825 271.625 195.895 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[3]

PIN DB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL2 ;
RECT 204.645 0.0 205.715 0.64 ;
LAYER METAL3 ;
RECT 204.645 0.0 205.715 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[3]

PIN QA[2]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 218.065 271.625 219.135 272.265 ;
LAYER METAL2 ;
RECT 218.065 271.625 219.135 272.265 ;
LAYER METAL3 ;
RECT 218.065 271.625 219.135 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[2]

PIN DB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL2 ;
RECT 227.885 0.0 228.955 0.64 ;
LAYER METAL3 ;
RECT 227.885 0.0 228.955 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[2]

PIN QA[1]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 241.305 271.625 242.375 272.265 ;
LAYER METAL2 ;
RECT 241.305 271.625 242.375 272.265 ;
LAYER METAL3 ;
RECT 241.305 271.625 242.375 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[1]

PIN DB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL2 ;
RECT 251.125 0.0 252.195 0.64 ;
LAYER METAL3 ;
RECT 251.125 0.0 252.195 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[1]

PIN QA[0]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 264.545 271.625 265.615 272.265 ;
LAYER METAL2 ;
RECT 264.545 271.625 265.615 272.265 ;
LAYER METAL3 ;
RECT 264.545 271.625 265.615 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[0]

PIN DB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL2 ;
RECT 274.365 0.0 275.435 0.64 ;
LAYER METAL3 ;
RECT 274.365 0.0 275.435 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[0]

PIN CLKB
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL2 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL3 ;
RECT 297.105 0.0 297.605 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKB

PIN AA[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 297.655 271.625 298.905 272.265 ;
LAYER METAL2 ;
RECT 297.655 271.625 298.905 272.265 ;
LAYER METAL3 ;
RECT 297.655 271.625 298.905 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[0]

PIN AA[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 302.505 271.625 303.755 272.265 ;
LAYER METAL2 ;
RECT 302.505 271.625 303.755 272.265 ;
LAYER METAL3 ;
RECT 302.505 271.625 303.755 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[1]

PIN CENB
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL2 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL3 ;
RECT 306.72 0.0 307.22 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENB

PIN AA[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 312.875 271.625 314.525 272.265 ;
LAYER METAL2 ;
RECT 312.875 271.625 314.125 272.265 ;
LAYER METAL3 ;
RECT 312.875 271.625 314.125 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[4]

PIN AA[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 320.815 271.625 322.465 272.265 ;
LAYER METAL2 ;
RECT 320.815 271.625 322.065 272.265 ;
LAYER METAL3 ;
RECT 320.815 271.625 322.065 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[3]

PIN AB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 323.45 0.0 325.015 0.64 ;
LAYER METAL2 ;
RECT 323.765 0.0 325.015 0.64 ;
LAYER METAL3 ;
RECT 323.765 0.0 325.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[8]

PIN AA[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.755 271.625 330.405 272.265 ;
LAYER METAL2 ;
RECT 328.755 271.625 330.005 272.265 ;
LAYER METAL3 ;
RECT 328.755 271.625 330.005 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[2]

PIN AB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 329.21 0.0 330.775 0.64 ;
LAYER METAL2 ;
RECT 329.525 0.0 330.775 0.64 ;
LAYER METAL3 ;
RECT 329.525 0.0 330.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[7]

PIN AA[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.365 271.625 335.93 272.265 ;
LAYER METAL2 ;
RECT 334.365 271.625 335.615 272.265 ;
LAYER METAL3 ;
RECT 334.365 271.625 335.615 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[5]

PIN AB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.97 0.0 336.535 0.64 ;
LAYER METAL2 ;
RECT 335.285 0.0 336.535 0.64 ;
LAYER METAL3 ;
RECT 335.285 0.0 336.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[6]

PIN AA[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.125 271.625 341.69 272.265 ;
LAYER METAL2 ;
RECT 340.125 271.625 341.375 272.265 ;
LAYER METAL3 ;
RECT 340.125 271.625 341.375 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[6]

PIN AB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.73 0.0 342.295 0.64 ;
LAYER METAL2 ;
RECT 341.045 0.0 342.295 0.64 ;
LAYER METAL3 ;
RECT 341.045 0.0 342.295 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[5]

PIN AA[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 345.885 271.625 347.45 272.265 ;
LAYER METAL2 ;
RECT 345.885 271.625 347.135 272.265 ;
LAYER METAL3 ;
RECT 345.885 271.625 347.135 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[7]

PIN AB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 346.255 0.0 347.905 0.64 ;
LAYER METAL2 ;
RECT 346.655 0.0 347.905 0.64 ;
LAYER METAL3 ;
RECT 346.655 0.0 347.905 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[2]

PIN AA[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 351.645 271.625 353.21 272.265 ;
LAYER METAL2 ;
RECT 351.645 271.625 352.895 272.265 ;
LAYER METAL3 ;
RECT 351.645 271.625 352.895 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[8]

PIN AB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 354.195 0.0 355.845 0.64 ;
LAYER METAL2 ;
RECT 354.595 0.0 355.845 0.64 ;
LAYER METAL3 ;
RECT 354.595 0.0 355.845 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[3]

PIN AB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 362.135 0.0 363.785 0.64 ;
LAYER METAL2 ;
RECT 362.535 0.0 363.785 0.64 ;
LAYER METAL3 ;
RECT 362.535 0.0 363.785 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[4]

PIN CENA
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 371.285 271.195 371.785 272.265 ;
LAYER METAL2 ;
RECT 371.285 271.195 371.785 272.265 ;
LAYER METAL3 ;
RECT 371.285 271.195 371.785 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENA

PIN AB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 372.905 0.0 374.155 0.64 ;
LAYER METAL2 ;
RECT 372.905 0.0 374.155 0.64 ;
LAYER METAL3 ;
RECT 372.905 0.0 374.155 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[1]

PIN AB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 377.755 0.0 379.005 0.64 ;
LAYER METAL2 ;
RECT 377.755 0.0 379.005 0.64 ;
LAYER METAL3 ;
RECT 377.755 0.0 379.005 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[0]

PIN CLKA
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 380.69 271.195 381.19 272.265 ;
LAYER METAL2 ;
RECT 380.69 271.195 381.19 272.265 ;
LAYER METAL3 ;
RECT 380.69 271.195 381.19 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKA

PIN DB[12]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 401.225 0.0 402.295 0.64 ;
LAYER METAL2 ;
RECT 401.225 0.0 402.295 0.64 ;
LAYER METAL3 ;
RECT 401.225 0.0 402.295 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[12]

PIN QA[12]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 411.045 271.625 412.115 272.265 ;
LAYER METAL2 ;
RECT 411.045 271.625 412.115 272.265 ;
LAYER METAL3 ;
RECT 411.045 271.625 412.115 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[12]

PIN DB[13]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 424.465 0.0 425.535 0.64 ;
LAYER METAL2 ;
RECT 424.465 0.0 425.535 0.64 ;
LAYER METAL3 ;
RECT 424.465 0.0 425.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[13]

PIN QA[13]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 434.285 271.625 435.355 272.265 ;
LAYER METAL2 ;
RECT 434.285 271.625 435.355 272.265 ;
LAYER METAL3 ;
RECT 434.285 271.625 435.355 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[13]

PIN DB[14]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 447.705 0.0 448.775 0.64 ;
LAYER METAL2 ;
RECT 447.705 0.0 448.775 0.64 ;
LAYER METAL3 ;
RECT 447.705 0.0 448.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[14]

PIN QA[14]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 457.525 271.625 458.595 272.265 ;
LAYER METAL2 ;
RECT 457.525 271.625 458.595 272.265 ;
LAYER METAL3 ;
RECT 457.525 271.625 458.595 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[14]

PIN DB[15]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 470.945 0.0 472.015 0.64 ;
LAYER METAL2 ;
RECT 470.945 0.0 472.015 0.64 ;
LAYER METAL3 ;
RECT 470.945 0.0 472.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[15]

PIN QA[15]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 480.765 271.625 481.835 272.265 ;
LAYER METAL2 ;
RECT 480.765 271.625 481.835 272.265 ;
LAYER METAL3 ;
RECT 480.765 271.625 481.835 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[15]

PIN DB[16]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 494.185 0.0 495.255 0.64 ;
LAYER METAL2 ;
RECT 494.185 0.0 495.255 0.64 ;
LAYER METAL3 ;
RECT 494.185 0.0 495.255 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[16]

PIN QA[16]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 504.005 271.625 505.075 272.265 ;
LAYER METAL2 ;
RECT 504.005 271.625 505.075 272.265 ;
LAYER METAL3 ;
RECT 504.005 271.625 505.075 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[16]

PIN DB[17]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 517.425 0.0 518.495 0.64 ;
LAYER METAL2 ;
RECT 517.425 0.0 518.495 0.64 ;
LAYER METAL3 ;
RECT 517.425 0.0 518.495 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[17]

PIN QA[17]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 527.245 271.625 528.315 272.265 ;
LAYER METAL2 ;
RECT 527.245 271.625 528.315 272.265 ;
LAYER METAL3 ;
RECT 527.245 271.625 528.315 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[17]

PIN DB[18]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 540.665 0.0 541.735 0.64 ;
LAYER METAL2 ;
RECT 540.665 0.0 541.735 0.64 ;
LAYER METAL3 ;
RECT 540.665 0.0 541.735 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[18]

PIN QA[18]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 550.485 271.625 551.555 272.265 ;
LAYER METAL2 ;
RECT 550.485 271.625 551.555 272.265 ;
LAYER METAL3 ;
RECT 550.485 271.625 551.555 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[18]

PIN DB[19]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 563.905 0.0 564.975 0.64 ;
LAYER METAL2 ;
RECT 563.905 0.0 564.975 0.64 ;
LAYER METAL3 ;
RECT 563.905 0.0 564.975 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[19]

PIN QA[19]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 573.725 271.625 574.795 272.265 ;
LAYER METAL2 ;
RECT 573.725 271.625 574.795 272.265 ;
LAYER METAL3 ;
RECT 573.725 271.625 574.795 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[19]

PIN DB[20]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 587.145 0.0 588.215 0.64 ;
LAYER METAL2 ;
RECT 587.145 0.0 588.215 0.64 ;
LAYER METAL3 ;
RECT 587.145 0.0 588.215 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[20]

PIN QA[20]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 596.965 271.625 598.035 272.265 ;
LAYER METAL2 ;
RECT 596.965 271.625 598.035 272.265 ;
LAYER METAL3 ;
RECT 596.965 271.625 598.035 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[20]

PIN DB[21]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 610.385 0.0 611.455 0.64 ;
LAYER METAL2 ;
RECT 610.385 0.0 611.455 0.64 ;
LAYER METAL3 ;
RECT 610.385 0.0 611.455 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[21]

PIN QA[21]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 620.205 271.625 621.275 272.265 ;
LAYER METAL2 ;
RECT 620.205 271.625 621.275 272.265 ;
LAYER METAL3 ;
RECT 620.205 271.625 621.275 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[21]

PIN DB[22]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 633.625 0.0 634.695 0.64 ;
LAYER METAL2 ;
RECT 633.625 0.0 634.695 0.64 ;
LAYER METAL3 ;
RECT 633.625 0.0 634.695 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[22]

PIN QA[22]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 643.445 271.625 644.515 272.265 ;
LAYER METAL2 ;
RECT 643.445 271.625 644.515 272.265 ;
LAYER METAL3 ;
RECT 643.445 271.625 644.515 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[22]

PIN DB[23]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 656.865 0.0 657.935 0.64 ;
LAYER METAL2 ;
RECT 656.865 0.0 657.935 0.64 ;
LAYER METAL3 ;
RECT 656.865 0.0 657.935 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[23]

PIN QA[23]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 666.685 271.625 667.755 272.265 ;
LAYER METAL2 ;
RECT 666.685 271.625 667.755 272.265 ;
LAYER METAL3 ;
RECT 666.685 271.625 667.755 272.265 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[23]

PIN VSS
DIRECTION INOUT ;
USE GROUND ;
PORT
LAYER METAL4 ;
RECT 279.475 0.0 283.475 272.265 ;
LAYER METAL4 ;
RECT 290.475 0.0 294.475 272.265 ;
LAYER METAL4 ;
RECT 301.475 0.0 305.475 272.265 ;
LAYER METAL4 ;
RECT 312.475 0.0 316.475 272.265 ;
LAYER METAL4 ;
RECT 323.475 0.0 327.475 272.265 ;
LAYER METAL4 ;
RECT 349.185 0.0 353.185 272.265 ;
LAYER METAL4 ;
RECT 360.185 0.0 364.185 272.265 ;
LAYER METAL4 ;
RECT 371.185 0.0 375.185 272.265 ;
LAYER METAL4 ;
RECT 382.185 0.0 386.185 272.265 ;
LAYER METAL4 ;
RECT 393.185 0.0 397.185 272.265 ;
LAYER METAL4 ;
RECT 267.855 0.0 271.855 272.265 ;
LAYER METAL4 ;
RECT 256.235 0.0 260.235 272.265 ;
LAYER METAL4 ;
RECT 244.615 0.0 248.615 272.265 ;
LAYER METAL4 ;
RECT 232.995 0.0 236.995 272.265 ;
LAYER METAL4 ;
RECT 221.375 0.0 225.375 272.265 ;
LAYER METAL4 ;
RECT 209.755 0.0 213.755 272.265 ;
LAYER METAL4 ;
RECT 198.135 0.0 202.135 272.265 ;
LAYER METAL4 ;
RECT 186.515 0.0 190.515 272.265 ;
LAYER METAL4 ;
RECT 174.895 0.0 178.895 272.265 ;
LAYER METAL4 ;
RECT 163.275 0.0 167.275 272.265 ;
LAYER METAL4 ;
RECT 151.655 0.0 155.655 272.265 ;
LAYER METAL4 ;
RECT 140.035 0.0 144.035 272.265 ;
LAYER METAL4 ;
RECT 128.415 0.0 132.415 272.265 ;
LAYER METAL4 ;
RECT 116.795 0.0 120.795 272.265 ;
LAYER METAL4 ;
RECT 105.175 0.0 109.175 272.265 ;
LAYER METAL4 ;
RECT 93.555 0.0 97.555 272.265 ;
LAYER METAL4 ;
RECT 81.935 0.0 85.935 272.265 ;
LAYER METAL4 ;
RECT 70.315 0.0 74.315 272.265 ;
LAYER METAL4 ;
RECT 58.695 0.0 62.695 272.265 ;
LAYER METAL4 ;
RECT 47.075 0.0 51.075 272.265 ;
LAYER METAL4 ;
RECT 35.455 0.0 39.455 272.265 ;
LAYER METAL4 ;
RECT 23.835 0.0 27.835 272.265 ;
LAYER METAL4 ;
RECT 12.215 0.0 16.215 272.265 ;
LAYER METAL4 ;
RECT 0.595 0.0 4.595 272.265 ;
LAYER METAL4 ;
RECT 404.805 0.0 408.805 272.265 ;
LAYER METAL4 ;
RECT 416.425 0.0 420.425 272.265 ;
LAYER METAL4 ;
RECT 428.045 0.0 432.045 272.265 ;
LAYER METAL4 ;
RECT 439.665 0.0 443.665 272.265 ;
LAYER METAL4 ;
RECT 451.285 0.0 455.285 272.265 ;
LAYER METAL4 ;
RECT 462.905 0.0 466.905 272.265 ;
LAYER METAL4 ;
RECT 474.525 0.0 478.525 272.265 ;
LAYER METAL4 ;
RECT 486.145 0.0 490.145 272.265 ;
LAYER METAL4 ;
RECT 497.765 0.0 501.765 272.265 ;
LAYER METAL4 ;
RECT 509.385 0.0 513.385 272.265 ;
LAYER METAL4 ;
RECT 521.005 0.0 525.005 272.265 ;
LAYER METAL4 ;
RECT 532.625 0.0 536.625 272.265 ;
LAYER METAL4 ;
RECT 544.245 0.0 548.245 272.265 ;
LAYER METAL4 ;
RECT 555.865 0.0 559.865 272.265 ;
LAYER METAL4 ;
RECT 567.485 0.0 571.485 272.265 ;
LAYER METAL4 ;
RECT 579.105 0.0 583.105 272.265 ;
LAYER METAL4 ;
RECT 590.725 0.0 594.725 272.265 ;
LAYER METAL4 ;
RECT 602.345 0.0 606.345 272.265 ;
LAYER METAL4 ;
RECT 613.965 0.0 617.965 272.265 ;
LAYER METAL4 ;
RECT 625.585 0.0 629.585 272.265 ;
LAYER METAL4 ;
RECT 637.205 0.0 641.205 272.265 ;
LAYER METAL4 ;
RECT 648.825 0.0 652.825 272.265 ;
LAYER METAL4 ;
RECT 660.445 0.0 664.445 272.265 ;
LAYER METAL4 ;
RECT 672.065 0.0 676.065 272.265 ;
END
END VSS

PIN VDD
DIRECTION INOUT ;
USE POWER ;
PORT
LAYER METAL4 ;
RECT 284.975 0.0 288.975 272.265 ;
LAYER METAL4 ;
RECT 295.975 0.0 299.975 272.265 ;
LAYER METAL4 ;
RECT 306.975 0.0 310.975 272.265 ;
LAYER METAL4 ;
RECT 317.975 0.0 321.975 272.265 ;
LAYER METAL4 ;
RECT 328.975 0.0 332.975 272.265 ;
LAYER METAL4 ;
RECT 343.685 0.0 347.685 272.265 ;
LAYER METAL4 ;
RECT 354.685 0.0 358.685 272.265 ;
LAYER METAL4 ;
RECT 365.685 0.0 369.685 272.265 ;
LAYER METAL4 ;
RECT 376.685 0.0 380.685 272.265 ;
LAYER METAL4 ;
RECT 387.685 0.0 391.685 272.265 ;
LAYER METAL4 ;
RECT 273.665 0.0 277.665 272.265 ;
LAYER METAL4 ;
RECT 262.045 0.0 266.045 272.265 ;
LAYER METAL4 ;
RECT 250.425 0.0 254.425 272.265 ;
LAYER METAL4 ;
RECT 238.805 0.0 242.805 272.265 ;
LAYER METAL4 ;
RECT 227.185 0.0 231.185 272.265 ;
LAYER METAL4 ;
RECT 215.565 0.0 219.565 272.265 ;
LAYER METAL4 ;
RECT 203.945 0.0 207.945 272.265 ;
LAYER METAL4 ;
RECT 192.325 0.0 196.325 272.265 ;
LAYER METAL4 ;
RECT 180.705 0.0 184.705 272.265 ;
LAYER METAL4 ;
RECT 169.085 0.0 173.085 272.265 ;
LAYER METAL4 ;
RECT 157.465 0.0 161.465 272.265 ;
LAYER METAL4 ;
RECT 145.845 0.0 149.845 272.265 ;
LAYER METAL4 ;
RECT 134.225 0.0 138.225 272.265 ;
LAYER METAL4 ;
RECT 122.605 0.0 126.605 272.265 ;
LAYER METAL4 ;
RECT 110.985 0.0 114.985 272.265 ;
LAYER METAL4 ;
RECT 99.365 0.0 103.365 272.265 ;
LAYER METAL4 ;
RECT 87.745 0.0 91.745 272.265 ;
LAYER METAL4 ;
RECT 76.125 0.0 80.125 272.265 ;
LAYER METAL4 ;
RECT 64.505 0.0 68.505 272.265 ;
LAYER METAL4 ;
RECT 52.885 0.0 56.885 272.265 ;
LAYER METAL4 ;
RECT 41.265 0.0 45.265 272.265 ;
LAYER METAL4 ;
RECT 29.645 0.0 33.645 272.265 ;
LAYER METAL4 ;
RECT 18.025 0.0 22.025 272.265 ;
LAYER METAL4 ;
RECT 6.405 0.0 10.405 272.265 ;
LAYER METAL4 ;
RECT 398.995 0.0 402.995 272.265 ;
LAYER METAL4 ;
RECT 410.615 0.0 414.615 272.265 ;
LAYER METAL4 ;
RECT 422.235 0.0 426.235 272.265 ;
LAYER METAL4 ;
RECT 433.855 0.0 437.855 272.265 ;
LAYER METAL4 ;
RECT 445.475 0.0 449.475 272.265 ;
LAYER METAL4 ;
RECT 457.095 0.0 461.095 272.265 ;
LAYER METAL4 ;
RECT 468.715 0.0 472.715 272.265 ;
LAYER METAL4 ;
RECT 480.335 0.0 484.335 272.265 ;
LAYER METAL4 ;
RECT 491.955 0.0 495.955 272.265 ;
LAYER METAL4 ;
RECT 503.575 0.0 507.575 272.265 ;
LAYER METAL4 ;
RECT 515.195 0.0 519.195 272.265 ;
LAYER METAL4 ;
RECT 526.815 0.0 530.815 272.265 ;
LAYER METAL4 ;
RECT 538.435 0.0 542.435 272.265 ;
LAYER METAL4 ;
RECT 550.055 0.0 554.055 272.265 ;
LAYER METAL4 ;
RECT 561.675 0.0 565.675 272.265 ;
LAYER METAL4 ;
RECT 573.295 0.0 577.295 272.265 ;
LAYER METAL4 ;
RECT 584.915 0.0 588.915 272.265 ;
LAYER METAL4 ;
RECT 596.535 0.0 600.535 272.265 ;
LAYER METAL4 ;
RECT 608.155 0.0 612.155 272.265 ;
LAYER METAL4 ;
RECT 619.775 0.0 623.775 272.265 ;
LAYER METAL4 ;
RECT 631.395 0.0 635.395 272.265 ;
LAYER METAL4 ;
RECT 643.015 0.0 647.015 272.265 ;
LAYER METAL4 ;
RECT 654.635 0.0 658.635 272.265 ;
LAYER METAL4 ;
RECT 666.255 0.0 670.255 272.265 ;
END
END VDD

OBS
LAYER VIA12 ;
RECT  0.000 0.000 676.660 272.265 ;
LAYER VIA23 ;
RECT  0.000 0.000 676.660 272.265 ;
LAYER VIA34 ;
RECT  0.000 0.000 676.660 272.265 ;
LAYER METAL1 ;
POLYGON 0.000 0.000 18.495 0.000 18.495 0.870 20.025 0.870 20.025 0.000
 41.735 0.000 41.735 0.870 43.265 0.870 43.265 0.000 64.975 0.000
 64.975 0.870 66.505 0.870 66.505 0.000 88.215 0.000 88.215 0.870
 89.745 0.870 89.745 0.000 111.455 0.000 111.455 0.870 112.985 0.870
 112.985 0.000 134.695 0.000 134.695 0.870 136.225 0.870 136.225 0.000
 157.935 0.000 157.935 0.870 159.465 0.870 159.465 0.000 181.175 0.000
 181.175 0.870 182.705 0.870 182.705 0.000 204.415 0.000 204.415 0.870
 205.945 0.870 205.945 0.000 227.655 0.000 227.655 0.870 229.185 0.870
 229.185 0.000 250.895 0.000 250.895 0.870 252.425 0.870 252.425 0.000
 274.135 0.000 274.135 0.870 275.665 0.870 275.665 0.000 296.875 0.000
 296.875 1.300 297.835 1.300 297.835 0.000 306.490 0.000 306.490 1.300
 307.450 1.300 307.450 0.000 323.220 0.000 323.220 0.870 325.245 0.870
 325.245 0.000 328.980 0.000 328.980 0.870 331.005 0.870 331.005 0.000
 334.740 0.000 334.740 0.870 336.765 0.870 336.765 0.000 340.500 0.000
 340.500 0.870 342.525 0.870 342.525 0.000 346.025 0.000 346.025 0.870
 348.135 0.870 348.135 0.000 353.965 0.000 353.965 0.870 356.075 0.870
 356.075 0.000 361.905 0.000 361.905 0.870 364.015 0.870 364.015 0.000
 372.675 0.000 372.675 0.870 374.385 0.870 374.385 0.000 377.525 0.000
 377.525 0.870 379.235 0.870 379.235 0.000 400.995 0.000 400.995 0.870
 402.525 0.870 402.525 0.000 424.235 0.000 424.235 0.870 425.765 0.870
 425.765 0.000 447.475 0.000 447.475 0.870 449.005 0.870 449.005 0.000
 470.715 0.000 470.715 0.870 472.245 0.870 472.245 0.000 493.955 0.000
 493.955 0.870 495.485 0.870 495.485 0.000 517.195 0.000 517.195 0.870
 518.725 0.870 518.725 0.000 540.435 0.000 540.435 0.870 541.965 0.870
 541.965 0.000 563.675 0.000 563.675 0.870 565.205 0.870 565.205 0.000
 586.915 0.000 586.915 0.870 588.445 0.870 588.445 0.000 610.155 0.000
 610.155 0.870 611.685 0.870 611.685 0.000 633.395 0.000 633.395 0.870
 634.925 0.870 634.925 0.000 656.635 0.000 656.635 0.870 658.165 0.870
 658.165 0.000 676.660 0.000 676.660 272.265 667.985 272.265 667.985 271.395 666.455 271.395 666.455 272.265
 644.745 272.265 644.745 271.395 643.215 271.395 643.215 272.265 621.505 272.265
 621.505 271.395 619.975 271.395 619.975 272.265 598.265 272.265 598.265 271.395
 596.735 271.395 596.735 272.265 575.025 272.265 575.025 271.395 573.495 271.395
 573.495 272.265 551.785 272.265 551.785 271.395 550.255 271.395 550.255 272.265
 528.545 272.265 528.545 271.395 527.015 271.395 527.015 272.265 505.305 272.265
 505.305 271.395 503.775 271.395 503.775 272.265 482.065 272.265 482.065 271.395
 480.535 271.395 480.535 272.265 458.825 272.265 458.825 271.395 457.295 271.395
 457.295 272.265 435.585 272.265 435.585 271.395 434.055 271.395 434.055 272.265
 412.345 272.265 412.345 271.395 410.815 271.395 410.815 272.265 381.420 272.265
 381.420 270.965 380.460 270.965 380.460 272.265 372.015 272.265 372.015 270.965
 371.055 270.965 371.055 272.265 353.440 272.265 353.440 271.395 351.415 271.395
 351.415 272.265 347.680 272.265 347.680 271.395 345.655 271.395 345.655 272.265
 341.920 272.265 341.920 271.395 339.895 271.395 339.895 272.265 336.160 272.265
 336.160 271.395 334.135 271.395 334.135 272.265 330.635 272.265 330.635 271.395
 328.525 271.395 328.525 272.265 322.695 272.265 322.695 271.395 320.585 271.395
 320.585 272.265 314.755 272.265 314.755 271.395 312.645 271.395 312.645 272.265
 303.985 272.265 303.985 271.395 302.275 271.395 302.275 272.265 299.135 272.265
 299.135 271.395 297.425 271.395 297.425 272.265 265.845 272.265 265.845 271.395
 264.315 271.395 264.315 272.265 242.605 272.265 242.605 271.395 241.075 271.395
 241.075 272.265 219.365 272.265 219.365 271.395 217.835 271.395 217.835 272.265
 196.125 272.265 196.125 271.395 194.595 271.395 194.595 272.265 172.885 272.265
 172.885 271.395 171.355 271.395 171.355 272.265 149.645 272.265 149.645 271.395
 148.115 271.395 148.115 272.265 126.405 272.265 126.405 271.395 124.875 271.395
 124.875 272.265 103.165 272.265 103.165 271.395 101.635 271.395 101.635 272.265
 79.925 272.265 79.925 271.395 78.395 271.395 78.395 272.265 56.685 272.265
 56.685 271.395 55.155 271.395 55.155 272.265 33.445 272.265 33.445 271.395
 31.915 271.395 31.915 272.265 10.205 272.265 10.205 271.395 8.675 271.395
 8.675 272.265 0.000 272.265 ;
LAYER METAL2 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 335.005 0.000 335.005 0.920 336.815 0.920 336.815 0.000 340.765 0.000
 340.765 0.920 342.575 0.920 342.575 0.000 346.375 0.000 346.375 0.920
 348.185 0.920 348.185 0.000 354.315 0.000 354.315 0.920 356.125 0.920
 356.125 0.000 362.255 0.000 362.255 0.920 364.065 0.920 364.065 0.000
 372.625 0.000 372.625 0.920 374.435 0.920 374.435 0.000 377.475 0.000
 377.475 0.920 379.285 0.920 379.285 0.000 400.945 0.000 400.945 0.920
 402.575 0.920 402.575 0.000 424.185 0.000 424.185 0.920 425.815 0.920
 425.815 0.000 447.425 0.000 447.425 0.920 449.055 0.920 449.055 0.000
 470.665 0.000 470.665 0.920 472.295 0.920 472.295 0.000 493.905 0.000
 493.905 0.920 495.535 0.920 495.535 0.000 517.145 0.000 517.145 0.920
 518.775 0.920 518.775 0.000 540.385 0.000 540.385 0.920 542.015 0.920
 542.015 0.000 563.625 0.000 563.625 0.920 565.255 0.920 565.255 0.000
 586.865 0.000 586.865 0.920 588.495 0.920 588.495 0.000 610.105 0.000
 610.105 0.920 611.735 0.920 611.735 0.000 633.345 0.000 633.345 0.920
 634.975 0.920 634.975 0.000 656.585 0.000 656.585 0.920 658.215 0.920
 658.215 0.000 676.660 0.000 676.660 272.265 668.035 272.265 668.035 271.345 666.405 271.345 666.405 272.265
 644.795 272.265 644.795 271.345 643.165 271.345 643.165 272.265 621.555 272.265
 621.555 271.345 619.925 271.345 619.925 272.265 598.315 272.265 598.315 271.345
 596.685 271.345 596.685 272.265 575.075 272.265 575.075 271.345 573.445 271.345
 573.445 272.265 551.835 272.265 551.835 271.345 550.205 271.345 550.205 272.265
 528.595 272.265 528.595 271.345 526.965 271.345 526.965 272.265 505.355 272.265
 505.355 271.345 503.725 271.345 503.725 272.265 482.115 272.265 482.115 271.345
 480.485 271.345 480.485 272.265 458.875 272.265 458.875 271.345 457.245 271.345
 457.245 272.265 435.635 272.265 435.635 271.345 434.005 271.345 434.005 272.265
 412.395 272.265 412.395 271.345 410.765 271.345 410.765 272.265 381.470 272.265
 381.470 270.915 380.410 270.915 380.410 272.265 372.065 272.265 372.065 270.915
 371.005 270.915 371.005 272.265 353.175 272.265 353.175 271.345 351.365 271.345
 351.365 272.265 347.415 272.265 347.415 271.345 345.605 271.345 345.605 272.265
 341.655 272.265 341.655 271.345 339.845 271.345 339.845 272.265 335.895 272.265
 335.895 271.345 334.085 271.345 334.085 272.265 330.285 272.265 330.285 271.345
 328.475 271.345 328.475 272.265 322.345 272.265 322.345 271.345 320.535 271.345
 320.535 272.265 314.405 272.265 314.405 271.345 312.595 271.345 312.595 272.265
 304.035 272.265 304.035 271.345 302.225 271.345 302.225 272.265 299.185 272.265
 299.185 271.345 297.375 271.345 297.375 272.265 265.895 272.265 265.895 271.345
 264.265 271.345 264.265 272.265 242.655 272.265 242.655 271.345 241.025 271.345
 241.025 272.265 219.415 272.265 219.415 271.345 217.785 271.345 217.785 272.265
 196.175 272.265 196.175 271.345 194.545 271.345 194.545 272.265 172.935 272.265
 172.935 271.345 171.305 271.345 171.305 272.265 149.695 272.265 149.695 271.345
 148.065 271.345 148.065 272.265 126.455 272.265 126.455 271.345 124.825 271.345
 124.825 272.265 103.215 272.265 103.215 271.345 101.585 271.345 101.585 272.265
 79.975 272.265 79.975 271.345 78.345 271.345 78.345 272.265 56.735 272.265
 56.735 271.345 55.105 271.345 55.105 272.265 33.495 272.265 33.495 271.345
 31.865 271.345 31.865 272.265 10.255 272.265 10.255 271.345 8.625 271.345
 8.625 272.265 0.000 272.265 ;
LAYER METAL3 ;
POLYGON 0.000 0.000 18.445 0.000 18.445 0.920 20.075 0.920 20.075 0.000
 41.685 0.000 41.685 0.920 43.315 0.920 43.315 0.000 64.925 0.000
 64.925 0.920 66.555 0.920 66.555 0.000 88.165 0.000 88.165 0.920
 89.795 0.920 89.795 0.000 111.405 0.000 111.405 0.920 113.035 0.920
 113.035 0.000 134.645 0.000 134.645 0.920 136.275 0.920 136.275 0.000
 157.885 0.000 157.885 0.920 159.515 0.920 159.515 0.000 181.125 0.000
 181.125 0.920 182.755 0.920 182.755 0.000 204.365 0.000 204.365 0.920
 205.995 0.920 205.995 0.000 227.605 0.000 227.605 0.920 229.235 0.920
 229.235 0.000 250.845 0.000 250.845 0.920 252.475 0.920 252.475 0.000
 274.085 0.000 274.085 0.920 275.715 0.920 275.715 0.000 296.825 0.000
 296.825 1.350 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350
 307.500 1.350 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920
 325.295 0.000 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000
 335.005 0.000 335.005 0.920 336.815 0.920 336.815 0.000 340.765 0.000
 340.765 0.920 342.575 0.920 342.575 0.000 346.375 0.000 346.375 0.920
 348.185 0.920 348.185 0.000 354.315 0.000 354.315 0.920 356.125 0.920
 356.125 0.000 362.255 0.000 362.255 0.920 364.065 0.920 364.065 0.000
 372.625 0.000 372.625 0.920 374.435 0.920 374.435 0.000 377.475 0.000
 377.475 0.920 379.285 0.920 379.285 0.000 400.945 0.000 400.945 0.920
 402.575 0.920 402.575 0.000 424.185 0.000 424.185 0.920 425.815 0.920
 425.815 0.000 447.425 0.000 447.425 0.920 449.055 0.920 449.055 0.000
 470.665 0.000 470.665 0.920 472.295 0.920 472.295 0.000 493.905 0.000
 493.905 0.920 495.535 0.920 495.535 0.000 517.145 0.000 517.145 0.920
 518.775 0.920 518.775 0.000 540.385 0.000 540.385 0.920 542.015 0.920
 542.015 0.000 563.625 0.000 563.625 0.920 565.255 0.920 565.255 0.000
 586.865 0.000 586.865 0.920 588.495 0.920 588.495 0.000 610.105 0.000
 610.105 0.920 611.735 0.920 611.735 0.000 633.345 0.000 633.345 0.920
 634.975 0.920 634.975 0.000 656.585 0.000 656.585 0.920 658.215 0.920
 658.215 0.000 676.660 0.000 676.660 272.265 668.035 272.265 668.035 271.345 666.405 271.345 666.405 272.265
 644.795 272.265 644.795 271.345 643.165 271.345 643.165 272.265 621.555 272.265
 621.555 271.345 619.925 271.345 619.925 272.265 598.315 272.265 598.315 271.345
 596.685 271.345 596.685 272.265 575.075 272.265 575.075 271.345 573.445 271.345
 573.445 272.265 551.835 272.265 551.835 271.345 550.205 271.345 550.205 272.265
 528.595 272.265 528.595 271.345 526.965 271.345 526.965 272.265 505.355 272.265
 505.355 271.345 503.725 271.345 503.725 272.265 482.115 272.265 482.115 271.345
 480.485 271.345 480.485 272.265 458.875 272.265 458.875 271.345 457.245 271.345
 457.245 272.265 435.635 272.265 435.635 271.345 434.005 271.345 434.005 272.265
 412.395 272.265 412.395 271.345 410.765 271.345 410.765 272.265 381.470 272.265
 381.470 270.915 380.410 270.915 380.410 272.265 372.065 272.265 372.065 270.915
 371.005 270.915 371.005 272.265 353.175 272.265 353.175 271.345 351.365 271.345
 351.365 272.265 347.415 272.265 347.415 271.345 345.605 271.345 345.605 272.265
 341.655 272.265 341.655 271.345 339.845 271.345 339.845 272.265 335.895 272.265
 335.895 271.345 334.085 271.345 334.085 272.265 330.285 272.265 330.285 271.345
 328.475 271.345 328.475 272.265 322.345 272.265 322.345 271.345 320.535 271.345
 320.535 272.265 314.405 272.265 314.405 271.345 312.595 271.345 312.595 272.265
 304.035 272.265 304.035 271.345 302.225 271.345 302.225 272.265 299.185 272.265
 299.185 271.345 297.375 271.345 297.375 272.265 265.895 272.265 265.895 271.345
 264.265 271.345 264.265 272.265 242.655 272.265 242.655 271.345 241.025 271.345
 241.025 272.265 219.415 272.265 219.415 271.345 217.785 271.345 217.785 272.265
 196.175 272.265 196.175 271.345 194.545 271.345 194.545 272.265 172.935 272.265
 172.935 271.345 171.305 271.345 171.305 272.265 149.695 272.265 149.695 271.345
 148.065 271.345 148.065 272.265 126.455 272.265 126.455 271.345 124.825 271.345
 124.825 272.265 103.215 272.265 103.215 271.345 101.585 271.345 101.585 272.265
 79.975 272.265 79.975 271.345 78.345 271.345 78.345 272.265 56.735 272.265
 56.735 271.345 55.105 271.345 55.105 272.265 33.495 272.265 33.495 271.345
 31.865 271.345 31.865 272.265 10.255 272.265 10.255 271.345 8.625 271.345
 8.625 272.265 0.000 272.265 ;
END
END RAM512
END LIBRARY
