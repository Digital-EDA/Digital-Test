#     Copyright (c) 2023 SMIC                                                       
#     Filename:      FRAM512.lef                                                   
#     IP code:       S018RF2P                                                         
#     Version:       0.2.b                                                        
#     CreateDate:    Wed May 31 22:21:50 CST 2023                                                     
                    
#    LEF for 2-PORT Register File                                                               
#    SMIC 0.18um G Logic Process                                                       
#    Configuration: -instname FRAM512 -rows 256 -bits 48 -mux 2  



# DISCLAIMER                                                                           #
#                                                                                      #  
#   SMIC hereby provides the quality information to you but makes no claims,           #
# promises or guarantees about the accuracy, completeness, or adequacy of the          #
# information herein. The information contained herein is provided on an "AS IS"       #
# basis without any warranty, and SMIC assumes no obligation to provide support        #
# of any kind or otherwise maintain the information.                                   #  
#   SMIC disclaims any representation that the information does not infringe any       #
# intellectual property rights or proprietary rights of any third parties. SMIC        #
# makes no other warranty, whether express, implied or statutory as to any             #
# matter whatsoever, including but not limited to the accuracy or sufficiency of       #
# any information or the merchantability and fitness for a particular purpose.         #
# Neither SMIC nor any of its representatives shall be liable for any cause of         #
# action incurred to connect to this service.                                          #  
#                                                                                      #
# STATEMENT OF USE AND CONFIDENTIALITY                                                 #  
#                                                                                      #  
#   The following/attached material contains confidential and proprietary              #  
# information of SMIC. This material is based upon information which SMIC              #  
# considers reliable, but SMIC neither represents nor warrants that such               #
# information is accurate or complete, and it must not be relied upon as such.         #
# This information was prepared for informational purposes and is for the use          #
# by SMIC's customer only. SMIC reserves the right to make changes in the              #  
# information at any time without notice.                                              #  
#   No part of this information may be reproduced, transmitted, transcribed,           #  
# stored in a retrieval system, or translated into any human or computer               # 
# language, in any form or by any means, electronic, mechanical, magnetic,             #  
# optical, chemical, manual, or otherwise, without the prior written consent of        #
# SMIC. Any unauthorized use or disclosure of this material is strictly                #  
# prohibited and may be unlawful. By accepting this material, the receiving            #  
# party shall be deemed to have acknowledged, accepted, and agreed to be bound         #
# by the foregoing limitations and restrictions. Thank you.                            #  
#                                                                                      #  


MACRO FRAM512
CLASS BLOCK ;
ORIGIN 0 0 ;
SIZE 676.66 BY 496.905 ;
SYMMETRY X Y R90 ;

PIN DB[23]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 2.825 0.0 3.895 0.64 ;
LAYER METAL2 ;
RECT 2.825 0.0 3.895 0.64 ;
LAYER METAL3 ;
RECT 2.825 0.0 3.895 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[23]

PIN QA[23]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 12.645 496.265 13.715 496.905 ;
LAYER METAL2 ;
RECT 12.645 496.265 13.715 496.905 ;
LAYER METAL3 ;
RECT 12.645 496.265 13.715 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[23]

PIN QA[22]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 14.715 496.265 15.785 496.905 ;
LAYER METAL2 ;
RECT 14.715 496.265 15.785 496.905 ;
LAYER METAL3 ;
RECT 14.715 496.265 15.785 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[22]

PIN DB[22]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 24.535 0.0 25.605 0.64 ;
LAYER METAL2 ;
RECT 24.535 0.0 25.605 0.64 ;
LAYER METAL3 ;
RECT 24.535 0.0 25.605 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[22]

PIN DB[21]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 26.065 0.0 27.135 0.64 ;
LAYER METAL2 ;
RECT 26.065 0.0 27.135 0.64 ;
LAYER METAL3 ;
RECT 26.065 0.0 27.135 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[21]

PIN QA[21]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 35.885 496.265 36.955 496.905 ;
LAYER METAL2 ;
RECT 35.885 496.265 36.955 496.905 ;
LAYER METAL3 ;
RECT 35.885 496.265 36.955 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[21]

PIN QA[20]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 37.955 496.265 39.025 496.905 ;
LAYER METAL2 ;
RECT 37.955 496.265 39.025 496.905 ;
LAYER METAL3 ;
RECT 37.955 496.265 39.025 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[20]

PIN DB[20]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 47.775 0.0 48.845 0.64 ;
LAYER METAL2 ;
RECT 47.775 0.0 48.845 0.64 ;
LAYER METAL3 ;
RECT 47.775 0.0 48.845 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[20]

PIN DB[19]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 49.305 0.0 50.375 0.64 ;
LAYER METAL2 ;
RECT 49.305 0.0 50.375 0.64 ;
LAYER METAL3 ;
RECT 49.305 0.0 50.375 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[19]

PIN QA[19]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 59.125 496.265 60.195 496.905 ;
LAYER METAL2 ;
RECT 59.125 496.265 60.195 496.905 ;
LAYER METAL3 ;
RECT 59.125 496.265 60.195 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[19]

PIN QA[18]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 61.195 496.265 62.265 496.905 ;
LAYER METAL2 ;
RECT 61.195 496.265 62.265 496.905 ;
LAYER METAL3 ;
RECT 61.195 496.265 62.265 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[18]

PIN DB[18]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 71.015 0.0 72.085 0.64 ;
LAYER METAL2 ;
RECT 71.015 0.0 72.085 0.64 ;
LAYER METAL3 ;
RECT 71.015 0.0 72.085 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[18]

PIN DB[17]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 72.545 0.0 73.615 0.64 ;
LAYER METAL2 ;
RECT 72.545 0.0 73.615 0.64 ;
LAYER METAL3 ;
RECT 72.545 0.0 73.615 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[17]

PIN QA[17]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 82.365 496.265 83.435 496.905 ;
LAYER METAL2 ;
RECT 82.365 496.265 83.435 496.905 ;
LAYER METAL3 ;
RECT 82.365 496.265 83.435 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[17]

PIN QA[16]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 84.435 496.265 85.505 496.905 ;
LAYER METAL2 ;
RECT 84.435 496.265 85.505 496.905 ;
LAYER METAL3 ;
RECT 84.435 496.265 85.505 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[16]

PIN DB[16]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 94.255 0.0 95.325 0.64 ;
LAYER METAL2 ;
RECT 94.255 0.0 95.325 0.64 ;
LAYER METAL3 ;
RECT 94.255 0.0 95.325 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[16]

PIN DB[15]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 95.785 0.0 96.855 0.64 ;
LAYER METAL2 ;
RECT 95.785 0.0 96.855 0.64 ;
LAYER METAL3 ;
RECT 95.785 0.0 96.855 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[15]

PIN QA[15]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 105.605 496.265 106.675 496.905 ;
LAYER METAL2 ;
RECT 105.605 496.265 106.675 496.905 ;
LAYER METAL3 ;
RECT 105.605 496.265 106.675 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[15]

PIN QA[14]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 107.675 496.265 108.745 496.905 ;
LAYER METAL2 ;
RECT 107.675 496.265 108.745 496.905 ;
LAYER METAL3 ;
RECT 107.675 496.265 108.745 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[14]

PIN DB[14]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 117.495 0.0 118.565 0.64 ;
LAYER METAL2 ;
RECT 117.495 0.0 118.565 0.64 ;
LAYER METAL3 ;
RECT 117.495 0.0 118.565 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[14]

PIN DB[13]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 119.025 0.0 120.095 0.64 ;
LAYER METAL2 ;
RECT 119.025 0.0 120.095 0.64 ;
LAYER METAL3 ;
RECT 119.025 0.0 120.095 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[13]

PIN QA[13]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 128.845 496.265 129.915 496.905 ;
LAYER METAL2 ;
RECT 128.845 496.265 129.915 496.905 ;
LAYER METAL3 ;
RECT 128.845 496.265 129.915 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[13]

PIN QA[12]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 130.915 496.265 131.985 496.905 ;
LAYER METAL2 ;
RECT 130.915 496.265 131.985 496.905 ;
LAYER METAL3 ;
RECT 130.915 496.265 131.985 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[12]

PIN DB[12]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 140.735 0.0 141.805 0.64 ;
LAYER METAL2 ;
RECT 140.735 0.0 141.805 0.64 ;
LAYER METAL3 ;
RECT 140.735 0.0 141.805 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[12]

PIN DB[11]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 142.265 0.0 143.335 0.64 ;
LAYER METAL2 ;
RECT 142.265 0.0 143.335 0.64 ;
LAYER METAL3 ;
RECT 142.265 0.0 143.335 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[11]

PIN QA[11]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 152.085 496.265 153.155 496.905 ;
LAYER METAL2 ;
RECT 152.085 496.265 153.155 496.905 ;
LAYER METAL3 ;
RECT 152.085 496.265 153.155 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[11]

PIN QA[10]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 154.155 496.265 155.225 496.905 ;
LAYER METAL2 ;
RECT 154.155 496.265 155.225 496.905 ;
LAYER METAL3 ;
RECT 154.155 496.265 155.225 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[10]

PIN DB[10]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 163.975 0.0 165.045 0.64 ;
LAYER METAL2 ;
RECT 163.975 0.0 165.045 0.64 ;
LAYER METAL3 ;
RECT 163.975 0.0 165.045 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[10]

PIN DB[9]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 165.505 0.0 166.575 0.64 ;
LAYER METAL2 ;
RECT 165.505 0.0 166.575 0.64 ;
LAYER METAL3 ;
RECT 165.505 0.0 166.575 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[9]

PIN QA[9]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 175.325 496.265 176.395 496.905 ;
LAYER METAL2 ;
RECT 175.325 496.265 176.395 496.905 ;
LAYER METAL3 ;
RECT 175.325 496.265 176.395 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[9]

PIN QA[8]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 177.395 496.265 178.465 496.905 ;
LAYER METAL2 ;
RECT 177.395 496.265 178.465 496.905 ;
LAYER METAL3 ;
RECT 177.395 496.265 178.465 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[8]

PIN DB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 187.215 0.0 188.285 0.64 ;
LAYER METAL2 ;
RECT 187.215 0.0 188.285 0.64 ;
LAYER METAL3 ;
RECT 187.215 0.0 188.285 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[8]

PIN DB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 188.745 0.0 189.815 0.64 ;
LAYER METAL2 ;
RECT 188.745 0.0 189.815 0.64 ;
LAYER METAL3 ;
RECT 188.745 0.0 189.815 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[7]

PIN QA[7]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 198.565 496.265 199.635 496.905 ;
LAYER METAL2 ;
RECT 198.565 496.265 199.635 496.905 ;
LAYER METAL3 ;
RECT 198.565 496.265 199.635 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[7]

PIN QA[6]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 200.635 496.265 201.705 496.905 ;
LAYER METAL2 ;
RECT 200.635 496.265 201.705 496.905 ;
LAYER METAL3 ;
RECT 200.635 496.265 201.705 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[6]

PIN DB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 210.455 0.0 211.525 0.64 ;
LAYER METAL2 ;
RECT 210.455 0.0 211.525 0.64 ;
LAYER METAL3 ;
RECT 210.455 0.0 211.525 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[6]

PIN DB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 211.985 0.0 213.055 0.64 ;
LAYER METAL2 ;
RECT 211.985 0.0 213.055 0.64 ;
LAYER METAL3 ;
RECT 211.985 0.0 213.055 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[5]

PIN QA[5]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 221.805 496.265 222.875 496.905 ;
LAYER METAL2 ;
RECT 221.805 496.265 222.875 496.905 ;
LAYER METAL3 ;
RECT 221.805 496.265 222.875 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[5]

PIN QA[4]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 223.875 496.265 224.945 496.905 ;
LAYER METAL2 ;
RECT 223.875 496.265 224.945 496.905 ;
LAYER METAL3 ;
RECT 223.875 496.265 224.945 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[4]

PIN DB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 233.695 0.0 234.765 0.64 ;
LAYER METAL2 ;
RECT 233.695 0.0 234.765 0.64 ;
LAYER METAL3 ;
RECT 233.695 0.0 234.765 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[4]

PIN DB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 235.225 0.0 236.295 0.64 ;
LAYER METAL2 ;
RECT 235.225 0.0 236.295 0.64 ;
LAYER METAL3 ;
RECT 235.225 0.0 236.295 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[3]

PIN QA[3]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 245.045 496.265 246.115 496.905 ;
LAYER METAL2 ;
RECT 245.045 496.265 246.115 496.905 ;
LAYER METAL3 ;
RECT 245.045 496.265 246.115 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[3]

PIN QA[2]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 247.115 496.265 248.185 496.905 ;
LAYER METAL2 ;
RECT 247.115 496.265 248.185 496.905 ;
LAYER METAL3 ;
RECT 247.115 496.265 248.185 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[2]

PIN DB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 256.935 0.0 258.005 0.64 ;
LAYER METAL2 ;
RECT 256.935 0.0 258.005 0.64 ;
LAYER METAL3 ;
RECT 256.935 0.0 258.005 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[2]

PIN DB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 258.465 0.0 259.535 0.64 ;
LAYER METAL2 ;
RECT 258.465 0.0 259.535 0.64 ;
LAYER METAL3 ;
RECT 258.465 0.0 259.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[1]

PIN QA[1]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 268.285 496.265 269.355 496.905 ;
LAYER METAL2 ;
RECT 268.285 496.265 269.355 496.905 ;
LAYER METAL3 ;
RECT 268.285 496.265 269.355 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[1]

PIN QA[0]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 270.355 496.265 271.425 496.905 ;
LAYER METAL2 ;
RECT 270.355 496.265 271.425 496.905 ;
LAYER METAL3 ;
RECT 270.355 496.265 271.425 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[0]

PIN DB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 280.175 0.0 281.245 0.64 ;
LAYER METAL2 ;
RECT 280.175 0.0 281.245 0.64 ;
LAYER METAL3 ;
RECT 280.175 0.0 281.245 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[0]

PIN CLKB
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL2 ;
RECT 297.105 0.0 297.605 1.07 ;
LAYER METAL3 ;
RECT 297.105 0.0 297.605 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKB

PIN AA[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 297.3 496.265 298.55 496.905 ;
LAYER METAL2 ;
RECT 297.3 496.265 298.55 496.905 ;
LAYER METAL3 ;
RECT 297.3 496.265 298.55 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[0]

PIN CENB
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL2 ;
RECT 306.72 0.0 307.22 1.07 ;
LAYER METAL3 ;
RECT 306.72 0.0 307.22 1.07 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENB

PIN AA[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 307.115 496.265 308.765 496.905 ;
LAYER METAL2 ;
RECT 307.115 496.265 308.365 496.905 ;
LAYER METAL3 ;
RECT 307.115 496.265 308.365 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[3]

PIN AA[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 315.055 496.265 316.705 496.905 ;
LAYER METAL2 ;
RECT 315.055 496.265 316.305 496.905 ;
LAYER METAL3 ;
RECT 315.055 496.265 316.305 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[2]

PIN AA[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 322.995 496.265 324.645 496.905 ;
LAYER METAL2 ;
RECT 322.995 496.265 324.245 496.905 ;
LAYER METAL3 ;
RECT 322.995 496.265 324.245 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[1]

PIN AB[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 323.45 0.0 325.015 0.64 ;
LAYER METAL2 ;
RECT 323.765 0.0 325.015 0.64 ;
LAYER METAL3 ;
RECT 323.765 0.0 325.015 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[8]

PIN AA[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 328.605 496.265 330.17 496.905 ;
LAYER METAL2 ;
RECT 328.605 496.265 329.855 496.905 ;
LAYER METAL3 ;
RECT 328.605 496.265 329.855 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[4]

PIN AB[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 329.21 0.0 330.775 0.64 ;
LAYER METAL2 ;
RECT 329.525 0.0 330.775 0.64 ;
LAYER METAL3 ;
RECT 329.525 0.0 330.775 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[7]

PIN AA[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.365 496.265 335.93 496.905 ;
LAYER METAL2 ;
RECT 334.365 496.265 335.615 496.905 ;
LAYER METAL3 ;
RECT 334.365 496.265 335.615 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[5]

PIN AB[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 334.97 0.0 336.535 0.64 ;
LAYER METAL2 ;
RECT 335.285 0.0 336.535 0.64 ;
LAYER METAL3 ;
RECT 335.285 0.0 336.535 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[6]

PIN AA[6]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.125 496.265 341.69 496.905 ;
LAYER METAL2 ;
RECT 340.125 496.265 341.375 496.905 ;
LAYER METAL3 ;
RECT 340.125 496.265 341.375 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[6]

PIN AB[5]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 340.73 0.0 342.295 0.64 ;
LAYER METAL2 ;
RECT 341.045 0.0 342.295 0.64 ;
LAYER METAL3 ;
RECT 341.045 0.0 342.295 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[5]

PIN AA[7]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 345.885 496.265 347.45 496.905 ;
LAYER METAL2 ;
RECT 345.885 496.265 347.135 496.905 ;
LAYER METAL3 ;
RECT 345.885 496.265 347.135 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[7]

PIN AB[4]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 346.49 0.0 348.055 0.64 ;
LAYER METAL2 ;
RECT 346.805 0.0 348.055 0.64 ;
LAYER METAL3 ;
RECT 346.805 0.0 348.055 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[4]

PIN AA[8]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 351.645 496.265 353.21 496.905 ;
LAYER METAL2 ;
RECT 351.645 496.265 352.895 496.905 ;
LAYER METAL3 ;
RECT 351.645 496.265 352.895 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AA[8]

PIN AB[1]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 352.015 0.0 353.665 0.64 ;
LAYER METAL2 ;
RECT 352.415 0.0 353.665 0.64 ;
LAYER METAL3 ;
RECT 352.415 0.0 353.665 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[1]

PIN AB[2]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 359.955 0.0 361.605 0.64 ;
LAYER METAL2 ;
RECT 360.355 0.0 361.605 0.64 ;
LAYER METAL3 ;
RECT 360.355 0.0 361.605 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[2]

PIN AB[3]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 367.895 0.0 369.545 0.64 ;
LAYER METAL2 ;
RECT 368.295 0.0 369.545 0.64 ;
LAYER METAL3 ;
RECT 368.295 0.0 369.545 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[3]

PIN CENA
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 371.285 495.835 371.785 496.905 ;
LAYER METAL2 ;
RECT 371.285 495.835 371.785 496.905 ;
LAYER METAL3 ;
RECT 371.285 495.835 371.785 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CENA

PIN AB[0]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 378.11 0.0 379.36 0.64 ;
LAYER METAL2 ;
RECT 378.11 0.0 379.36 0.64 ;
LAYER METAL3 ;
RECT 378.11 0.0 379.36 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END AB[0]

PIN CLKA
DIRECTION INPUT ;
USE CLOCK ;
PORT
LAYER METAL1 ;
RECT 380.69 495.835 381.19 496.905 ;
LAYER METAL2 ;
RECT 380.69 495.835 381.19 496.905 ;
LAYER METAL3 ;
RECT 380.69 495.835 381.19 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END CLKA

PIN DB[24]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 395.415 0.0 396.485 0.64 ;
LAYER METAL2 ;
RECT 395.415 0.0 396.485 0.64 ;
LAYER METAL3 ;
RECT 395.415 0.0 396.485 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[24]

PIN QA[24]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 405.235 496.265 406.305 496.905 ;
LAYER METAL2 ;
RECT 405.235 496.265 406.305 496.905 ;
LAYER METAL3 ;
RECT 405.235 496.265 406.305 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[24]

PIN QA[25]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 407.305 496.265 408.375 496.905 ;
LAYER METAL2 ;
RECT 407.305 496.265 408.375 496.905 ;
LAYER METAL3 ;
RECT 407.305 496.265 408.375 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[25]

PIN DB[25]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 417.125 0.0 418.195 0.64 ;
LAYER METAL2 ;
RECT 417.125 0.0 418.195 0.64 ;
LAYER METAL3 ;
RECT 417.125 0.0 418.195 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[25]

PIN DB[26]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 418.655 0.0 419.725 0.64 ;
LAYER METAL2 ;
RECT 418.655 0.0 419.725 0.64 ;
LAYER METAL3 ;
RECT 418.655 0.0 419.725 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[26]

PIN QA[26]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 428.475 496.265 429.545 496.905 ;
LAYER METAL2 ;
RECT 428.475 496.265 429.545 496.905 ;
LAYER METAL3 ;
RECT 428.475 496.265 429.545 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[26]

PIN QA[27]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 430.545 496.265 431.615 496.905 ;
LAYER METAL2 ;
RECT 430.545 496.265 431.615 496.905 ;
LAYER METAL3 ;
RECT 430.545 496.265 431.615 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[27]

PIN DB[27]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 440.365 0.0 441.435 0.64 ;
LAYER METAL2 ;
RECT 440.365 0.0 441.435 0.64 ;
LAYER METAL3 ;
RECT 440.365 0.0 441.435 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[27]

PIN DB[28]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 441.895 0.0 442.965 0.64 ;
LAYER METAL2 ;
RECT 441.895 0.0 442.965 0.64 ;
LAYER METAL3 ;
RECT 441.895 0.0 442.965 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[28]

PIN QA[28]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 451.715 496.265 452.785 496.905 ;
LAYER METAL2 ;
RECT 451.715 496.265 452.785 496.905 ;
LAYER METAL3 ;
RECT 451.715 496.265 452.785 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[28]

PIN QA[29]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 453.785 496.265 454.855 496.905 ;
LAYER METAL2 ;
RECT 453.785 496.265 454.855 496.905 ;
LAYER METAL3 ;
RECT 453.785 496.265 454.855 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[29]

PIN DB[29]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 463.605 0.0 464.675 0.64 ;
LAYER METAL2 ;
RECT 463.605 0.0 464.675 0.64 ;
LAYER METAL3 ;
RECT 463.605 0.0 464.675 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[29]

PIN DB[30]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 465.135 0.0 466.205 0.64 ;
LAYER METAL2 ;
RECT 465.135 0.0 466.205 0.64 ;
LAYER METAL3 ;
RECT 465.135 0.0 466.205 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[30]

PIN QA[30]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 474.955 496.265 476.025 496.905 ;
LAYER METAL2 ;
RECT 474.955 496.265 476.025 496.905 ;
LAYER METAL3 ;
RECT 474.955 496.265 476.025 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[30]

PIN QA[31]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 477.025 496.265 478.095 496.905 ;
LAYER METAL2 ;
RECT 477.025 496.265 478.095 496.905 ;
LAYER METAL3 ;
RECT 477.025 496.265 478.095 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[31]

PIN DB[31]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 486.845 0.0 487.915 0.64 ;
LAYER METAL2 ;
RECT 486.845 0.0 487.915 0.64 ;
LAYER METAL3 ;
RECT 486.845 0.0 487.915 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[31]

PIN DB[32]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 488.375 0.0 489.445 0.64 ;
LAYER METAL2 ;
RECT 488.375 0.0 489.445 0.64 ;
LAYER METAL3 ;
RECT 488.375 0.0 489.445 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[32]

PIN QA[32]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 498.195 496.265 499.265 496.905 ;
LAYER METAL2 ;
RECT 498.195 496.265 499.265 496.905 ;
LAYER METAL3 ;
RECT 498.195 496.265 499.265 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[32]

PIN QA[33]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 500.265 496.265 501.335 496.905 ;
LAYER METAL2 ;
RECT 500.265 496.265 501.335 496.905 ;
LAYER METAL3 ;
RECT 500.265 496.265 501.335 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[33]

PIN DB[33]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 510.085 0.0 511.155 0.64 ;
LAYER METAL2 ;
RECT 510.085 0.0 511.155 0.64 ;
LAYER METAL3 ;
RECT 510.085 0.0 511.155 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[33]

PIN DB[34]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 511.615 0.0 512.685 0.64 ;
LAYER METAL2 ;
RECT 511.615 0.0 512.685 0.64 ;
LAYER METAL3 ;
RECT 511.615 0.0 512.685 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[34]

PIN QA[34]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 521.435 496.265 522.505 496.905 ;
LAYER METAL2 ;
RECT 521.435 496.265 522.505 496.905 ;
LAYER METAL3 ;
RECT 521.435 496.265 522.505 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[34]

PIN QA[35]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 523.505 496.265 524.575 496.905 ;
LAYER METAL2 ;
RECT 523.505 496.265 524.575 496.905 ;
LAYER METAL3 ;
RECT 523.505 496.265 524.575 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[35]

PIN DB[35]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 533.325 0.0 534.395 0.64 ;
LAYER METAL2 ;
RECT 533.325 0.0 534.395 0.64 ;
LAYER METAL3 ;
RECT 533.325 0.0 534.395 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[35]

PIN DB[36]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 534.855 0.0 535.925 0.64 ;
LAYER METAL2 ;
RECT 534.855 0.0 535.925 0.64 ;
LAYER METAL3 ;
RECT 534.855 0.0 535.925 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[36]

PIN QA[36]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 544.675 496.265 545.745 496.905 ;
LAYER METAL2 ;
RECT 544.675 496.265 545.745 496.905 ;
LAYER METAL3 ;
RECT 544.675 496.265 545.745 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[36]

PIN QA[37]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 546.745 496.265 547.815 496.905 ;
LAYER METAL2 ;
RECT 546.745 496.265 547.815 496.905 ;
LAYER METAL3 ;
RECT 546.745 496.265 547.815 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[37]

PIN DB[37]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 556.565 0.0 557.635 0.64 ;
LAYER METAL2 ;
RECT 556.565 0.0 557.635 0.64 ;
LAYER METAL3 ;
RECT 556.565 0.0 557.635 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[37]

PIN DB[38]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 558.095 0.0 559.165 0.64 ;
LAYER METAL2 ;
RECT 558.095 0.0 559.165 0.64 ;
LAYER METAL3 ;
RECT 558.095 0.0 559.165 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[38]

PIN QA[38]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 567.915 496.265 568.985 496.905 ;
LAYER METAL2 ;
RECT 567.915 496.265 568.985 496.905 ;
LAYER METAL3 ;
RECT 567.915 496.265 568.985 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[38]

PIN QA[39]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 569.985 496.265 571.055 496.905 ;
LAYER METAL2 ;
RECT 569.985 496.265 571.055 496.905 ;
LAYER METAL3 ;
RECT 569.985 496.265 571.055 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[39]

PIN DB[39]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 579.805 0.0 580.875 0.64 ;
LAYER METAL2 ;
RECT 579.805 0.0 580.875 0.64 ;
LAYER METAL3 ;
RECT 579.805 0.0 580.875 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[39]

PIN DB[40]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 581.335 0.0 582.405 0.64 ;
LAYER METAL2 ;
RECT 581.335 0.0 582.405 0.64 ;
LAYER METAL3 ;
RECT 581.335 0.0 582.405 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[40]

PIN QA[40]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 591.155 496.265 592.225 496.905 ;
LAYER METAL2 ;
RECT 591.155 496.265 592.225 496.905 ;
LAYER METAL3 ;
RECT 591.155 496.265 592.225 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[40]

PIN QA[41]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 593.225 496.265 594.295 496.905 ;
LAYER METAL2 ;
RECT 593.225 496.265 594.295 496.905 ;
LAYER METAL3 ;
RECT 593.225 496.265 594.295 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[41]

PIN DB[41]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 603.045 0.0 604.115 0.64 ;
LAYER METAL2 ;
RECT 603.045 0.0 604.115 0.64 ;
LAYER METAL3 ;
RECT 603.045 0.0 604.115 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[41]

PIN DB[42]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 604.575 0.0 605.645 0.64 ;
LAYER METAL2 ;
RECT 604.575 0.0 605.645 0.64 ;
LAYER METAL3 ;
RECT 604.575 0.0 605.645 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[42]

PIN QA[42]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 614.395 496.265 615.465 496.905 ;
LAYER METAL2 ;
RECT 614.395 496.265 615.465 496.905 ;
LAYER METAL3 ;
RECT 614.395 496.265 615.465 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[42]

PIN QA[43]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 616.465 496.265 617.535 496.905 ;
LAYER METAL2 ;
RECT 616.465 496.265 617.535 496.905 ;
LAYER METAL3 ;
RECT 616.465 496.265 617.535 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[43]

PIN DB[43]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 626.285 0.0 627.355 0.64 ;
LAYER METAL2 ;
RECT 626.285 0.0 627.355 0.64 ;
LAYER METAL3 ;
RECT 626.285 0.0 627.355 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[43]

PIN DB[44]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 627.815 0.0 628.885 0.64 ;
LAYER METAL2 ;
RECT 627.815 0.0 628.885 0.64 ;
LAYER METAL3 ;
RECT 627.815 0.0 628.885 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[44]

PIN QA[44]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 637.635 496.265 638.705 496.905 ;
LAYER METAL2 ;
RECT 637.635 496.265 638.705 496.905 ;
LAYER METAL3 ;
RECT 637.635 496.265 638.705 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[44]

PIN QA[45]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 639.705 496.265 640.775 496.905 ;
LAYER METAL2 ;
RECT 639.705 496.265 640.775 496.905 ;
LAYER METAL3 ;
RECT 639.705 496.265 640.775 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[45]

PIN DB[45]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 649.525 0.0 650.595 0.64 ;
LAYER METAL2 ;
RECT 649.525 0.0 650.595 0.64 ;
LAYER METAL3 ;
RECT 649.525 0.0 650.595 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[45]

PIN DB[46]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 651.055 0.0 652.125 0.64 ;
LAYER METAL2 ;
RECT 651.055 0.0 652.125 0.64 ;
LAYER METAL3 ;
RECT 651.055 0.0 652.125 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[46]

PIN QA[46]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 660.875 496.265 661.945 496.905 ;
LAYER METAL2 ;
RECT 660.875 496.265 661.945 496.905 ;
LAYER METAL3 ;
RECT 660.875 496.265 661.945 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[46]

PIN QA[47]
DIRECTION OUTPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 662.945 496.265 664.015 496.905 ;
LAYER METAL2 ;
RECT 662.945 496.265 664.015 496.905 ;
LAYER METAL3 ;
RECT 662.945 496.265 664.015 496.905 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END QA[47]

PIN DB[47]
DIRECTION INPUT ;
USE SIGNAL ;
PORT
LAYER METAL1 ;
RECT 672.765 0.0 673.835 0.64 ;
LAYER METAL2 ;
RECT 672.765 0.0 673.835 0.64 ;
LAYER METAL3 ;
RECT 672.765 0.0 673.835 0.64 ;
END
ANTENNAGATEAREA 0.079 ;
ANTENNADIFFAREA 0.3738 ;
END DB[47]

PIN VSS
DIRECTION INOUT ;
USE GROUND ;
PORT
LAYER METAL4 ;
RECT 279.475 0.0 283.475 496.905 ;
LAYER METAL4 ;
RECT 290.475 0.0 294.475 496.905 ;
LAYER METAL4 ;
RECT 301.475 0.0 305.475 496.905 ;
LAYER METAL4 ;
RECT 312.475 0.0 316.475 496.905 ;
LAYER METAL4 ;
RECT 323.475 0.0 327.475 496.905 ;
LAYER METAL4 ;
RECT 349.185 0.0 353.185 496.905 ;
LAYER METAL4 ;
RECT 360.185 0.0 364.185 496.905 ;
LAYER METAL4 ;
RECT 371.185 0.0 375.185 496.905 ;
LAYER METAL4 ;
RECT 382.185 0.0 386.185 496.905 ;
LAYER METAL4 ;
RECT 393.185 0.0 397.185 496.905 ;
LAYER METAL4 ;
RECT 267.855 0.0 271.855 496.905 ;
LAYER METAL4 ;
RECT 256.235 0.0 260.235 496.905 ;
LAYER METAL4 ;
RECT 244.615 0.0 248.615 496.905 ;
LAYER METAL4 ;
RECT 232.995 0.0 236.995 496.905 ;
LAYER METAL4 ;
RECT 221.375 0.0 225.375 496.905 ;
LAYER METAL4 ;
RECT 209.755 0.0 213.755 496.905 ;
LAYER METAL4 ;
RECT 198.135 0.0 202.135 496.905 ;
LAYER METAL4 ;
RECT 186.515 0.0 190.515 496.905 ;
LAYER METAL4 ;
RECT 174.895 0.0 178.895 496.905 ;
LAYER METAL4 ;
RECT 163.275 0.0 167.275 496.905 ;
LAYER METAL4 ;
RECT 151.655 0.0 155.655 496.905 ;
LAYER METAL4 ;
RECT 140.035 0.0 144.035 496.905 ;
LAYER METAL4 ;
RECT 128.415 0.0 132.415 496.905 ;
LAYER METAL4 ;
RECT 116.795 0.0 120.795 496.905 ;
LAYER METAL4 ;
RECT 105.175 0.0 109.175 496.905 ;
LAYER METAL4 ;
RECT 93.555 0.0 97.555 496.905 ;
LAYER METAL4 ;
RECT 81.935 0.0 85.935 496.905 ;
LAYER METAL4 ;
RECT 70.315 0.0 74.315 496.905 ;
LAYER METAL4 ;
RECT 58.695 0.0 62.695 496.905 ;
LAYER METAL4 ;
RECT 47.075 0.0 51.075 496.905 ;
LAYER METAL4 ;
RECT 35.455 0.0 39.455 496.905 ;
LAYER METAL4 ;
RECT 23.835 0.0 27.835 496.905 ;
LAYER METAL4 ;
RECT 12.215 0.0 16.215 496.905 ;
LAYER METAL4 ;
RECT 0.595 0.0 4.595 496.905 ;
LAYER METAL4 ;
RECT 404.805 0.0 408.805 496.905 ;
LAYER METAL4 ;
RECT 416.425 0.0 420.425 496.905 ;
LAYER METAL4 ;
RECT 428.045 0.0 432.045 496.905 ;
LAYER METAL4 ;
RECT 439.665 0.0 443.665 496.905 ;
LAYER METAL4 ;
RECT 451.285 0.0 455.285 496.905 ;
LAYER METAL4 ;
RECT 462.905 0.0 466.905 496.905 ;
LAYER METAL4 ;
RECT 474.525 0.0 478.525 496.905 ;
LAYER METAL4 ;
RECT 486.145 0.0 490.145 496.905 ;
LAYER METAL4 ;
RECT 497.765 0.0 501.765 496.905 ;
LAYER METAL4 ;
RECT 509.385 0.0 513.385 496.905 ;
LAYER METAL4 ;
RECT 521.005 0.0 525.005 496.905 ;
LAYER METAL4 ;
RECT 532.625 0.0 536.625 496.905 ;
LAYER METAL4 ;
RECT 544.245 0.0 548.245 496.905 ;
LAYER METAL4 ;
RECT 555.865 0.0 559.865 496.905 ;
LAYER METAL4 ;
RECT 567.485 0.0 571.485 496.905 ;
LAYER METAL4 ;
RECT 579.105 0.0 583.105 496.905 ;
LAYER METAL4 ;
RECT 590.725 0.0 594.725 496.905 ;
LAYER METAL4 ;
RECT 602.345 0.0 606.345 496.905 ;
LAYER METAL4 ;
RECT 613.965 0.0 617.965 496.905 ;
LAYER METAL4 ;
RECT 625.585 0.0 629.585 496.905 ;
LAYER METAL4 ;
RECT 637.205 0.0 641.205 496.905 ;
LAYER METAL4 ;
RECT 648.825 0.0 652.825 496.905 ;
LAYER METAL4 ;
RECT 660.445 0.0 664.445 496.905 ;
LAYER METAL4 ;
RECT 672.065 0.0 676.065 496.905 ;
END
END VSS

PIN VDD
DIRECTION INOUT ;
USE POWER ;
PORT
LAYER METAL4 ;
RECT 284.975 0.0 288.975 496.905 ;
LAYER METAL4 ;
RECT 295.975 0.0 299.975 496.905 ;
LAYER METAL4 ;
RECT 306.975 0.0 310.975 496.905 ;
LAYER METAL4 ;
RECT 317.975 0.0 321.975 496.905 ;
LAYER METAL4 ;
RECT 328.975 0.0 332.975 496.905 ;
LAYER METAL4 ;
RECT 343.685 0.0 347.685 496.905 ;
LAYER METAL4 ;
RECT 354.685 0.0 358.685 496.905 ;
LAYER METAL4 ;
RECT 365.685 0.0 369.685 496.905 ;
LAYER METAL4 ;
RECT 376.685 0.0 380.685 496.905 ;
LAYER METAL4 ;
RECT 387.685 0.0 391.685 496.905 ;
LAYER METAL4 ;
RECT 273.665 0.0 277.665 496.905 ;
LAYER METAL4 ;
RECT 262.045 0.0 266.045 496.905 ;
LAYER METAL4 ;
RECT 250.425 0.0 254.425 496.905 ;
LAYER METAL4 ;
RECT 238.805 0.0 242.805 496.905 ;
LAYER METAL4 ;
RECT 227.185 0.0 231.185 496.905 ;
LAYER METAL4 ;
RECT 215.565 0.0 219.565 496.905 ;
LAYER METAL4 ;
RECT 203.945 0.0 207.945 496.905 ;
LAYER METAL4 ;
RECT 192.325 0.0 196.325 496.905 ;
LAYER METAL4 ;
RECT 180.705 0.0 184.705 496.905 ;
LAYER METAL4 ;
RECT 169.085 0.0 173.085 496.905 ;
LAYER METAL4 ;
RECT 157.465 0.0 161.465 496.905 ;
LAYER METAL4 ;
RECT 145.845 0.0 149.845 496.905 ;
LAYER METAL4 ;
RECT 134.225 0.0 138.225 496.905 ;
LAYER METAL4 ;
RECT 122.605 0.0 126.605 496.905 ;
LAYER METAL4 ;
RECT 110.985 0.0 114.985 496.905 ;
LAYER METAL4 ;
RECT 99.365 0.0 103.365 496.905 ;
LAYER METAL4 ;
RECT 87.745 0.0 91.745 496.905 ;
LAYER METAL4 ;
RECT 76.125 0.0 80.125 496.905 ;
LAYER METAL4 ;
RECT 64.505 0.0 68.505 496.905 ;
LAYER METAL4 ;
RECT 52.885 0.0 56.885 496.905 ;
LAYER METAL4 ;
RECT 41.265 0.0 45.265 496.905 ;
LAYER METAL4 ;
RECT 29.645 0.0 33.645 496.905 ;
LAYER METAL4 ;
RECT 18.025 0.0 22.025 496.905 ;
LAYER METAL4 ;
RECT 6.405 0.0 10.405 496.905 ;
LAYER METAL4 ;
RECT 398.995 0.0 402.995 496.905 ;
LAYER METAL4 ;
RECT 410.615 0.0 414.615 496.905 ;
LAYER METAL4 ;
RECT 422.235 0.0 426.235 496.905 ;
LAYER METAL4 ;
RECT 433.855 0.0 437.855 496.905 ;
LAYER METAL4 ;
RECT 445.475 0.0 449.475 496.905 ;
LAYER METAL4 ;
RECT 457.095 0.0 461.095 496.905 ;
LAYER METAL4 ;
RECT 468.715 0.0 472.715 496.905 ;
LAYER METAL4 ;
RECT 480.335 0.0 484.335 496.905 ;
LAYER METAL4 ;
RECT 491.955 0.0 495.955 496.905 ;
LAYER METAL4 ;
RECT 503.575 0.0 507.575 496.905 ;
LAYER METAL4 ;
RECT 515.195 0.0 519.195 496.905 ;
LAYER METAL4 ;
RECT 526.815 0.0 530.815 496.905 ;
LAYER METAL4 ;
RECT 538.435 0.0 542.435 496.905 ;
LAYER METAL4 ;
RECT 550.055 0.0 554.055 496.905 ;
LAYER METAL4 ;
RECT 561.675 0.0 565.675 496.905 ;
LAYER METAL4 ;
RECT 573.295 0.0 577.295 496.905 ;
LAYER METAL4 ;
RECT 584.915 0.0 588.915 496.905 ;
LAYER METAL4 ;
RECT 596.535 0.0 600.535 496.905 ;
LAYER METAL4 ;
RECT 608.155 0.0 612.155 496.905 ;
LAYER METAL4 ;
RECT 619.775 0.0 623.775 496.905 ;
LAYER METAL4 ;
RECT 631.395 0.0 635.395 496.905 ;
LAYER METAL4 ;
RECT 643.015 0.0 647.015 496.905 ;
LAYER METAL4 ;
RECT 654.635 0.0 658.635 496.905 ;
LAYER METAL4 ;
RECT 666.255 0.0 670.255 496.905 ;
END
END VDD

OBS
LAYER VIA12 ;
RECT  0.000 0.000 676.660 496.905 ;
LAYER VIA23 ;
RECT  0.000 0.000 676.660 496.905 ;
LAYER VIA34 ;
RECT  0.000 0.000 676.660 496.905 ;
LAYER METAL1 ;
POLYGON 0.000 0.000 2.595 0.000 2.595 0.870 4.125 0.870 4.125 0.000
 24.305 0.000 24.305 0.870 27.365 0.870 27.365 0.000 47.545 0.000
 47.545 0.870 49.075 0.870 49.075 0.000 49.075 0.000 49.075 0.870
 50.605 0.870 50.605 0.000 70.785 0.000 70.785 0.870 73.845 0.870
 73.845 0.000 94.025 0.000 94.025 0.870 97.085 0.870 97.085 0.000
 117.265 0.000 117.265 0.870 120.325 0.870 120.325 0.000 140.505 0.000
 140.505 0.870 143.565 0.870 143.565 0.000 163.745 0.000 163.745 0.870
 165.275 0.870 165.275 0.000 165.275 0.000 165.275 0.870 166.805 0.870
 166.805 0.000 186.985 0.000 186.985 0.870 188.515 0.870 188.515 0.000
 188.515 0.000 188.515 0.870 190.045 0.870 190.045 0.000 210.225 0.000
 210.225 0.870 211.755 0.870 211.755 0.000 211.755 0.000 211.755 0.870
 213.285 0.870 213.285 0.000 233.465 0.000 233.465 0.870 234.995 0.870
 234.995 0.000 234.995 0.000 234.995 0.870 236.525 0.870 236.525 0.000
 256.705 0.000 256.705 0.870 259.765 0.870 259.765 0.000 279.945 0.000
 279.945 0.870 281.475 0.870 281.475 0.000 296.875 0.000 296.875 1.300
 297.835 1.300 297.835 0.000 306.490 0.000 306.490 1.300 307.450 1.300
 307.450 0.000 323.220 0.000 323.220 0.870 325.245 0.870 325.245 0.000
 328.980 0.000 328.980 0.870 331.005 0.870 331.005 0.000 334.740 0.000
 334.740 0.870 336.765 0.870 336.765 0.000 340.500 0.000 340.500 0.870
 342.525 0.870 342.525 0.000 346.260 0.000 346.260 0.870 348.285 0.870
 348.285 0.000 351.785 0.000 351.785 0.870 353.895 0.870 353.895 0.000
 359.725 0.000 359.725 0.870 361.835 0.870 361.835 0.000 367.665 0.000
 367.665 0.870 369.775 0.870 369.775 0.000 377.880 0.000 377.880 0.870
 379.590 0.870 379.590 0.000 395.185 0.000 395.185 0.870 396.715 0.870
 396.715 0.000 416.895 0.000 416.895 0.870 419.955 0.870 419.955 0.000
 440.135 0.000 440.135 0.870 443.195 0.870 443.195 0.000 463.375 0.000
 463.375 0.870 466.435 0.870 466.435 0.000 486.615 0.000 486.615 0.870
 489.675 0.870 489.675 0.000 509.855 0.000 509.855 0.870 512.915 0.870
 512.915 0.000 533.095 0.000 533.095 0.870 536.155 0.870 536.155 0.000
 556.335 0.000 556.335 0.870 559.395 0.870 559.395 0.000 579.575 0.000
 579.575 0.870 582.635 0.870 582.635 0.000 602.815 0.000 602.815 0.870
 605.875 0.870 605.875 0.000 626.055 0.000 626.055 0.870 629.115 0.870
 629.115 0.000 649.295 0.000 649.295 0.870 652.355 0.870 652.355 0.000
 672.535 0.000 672.535 0.870 674.065 0.870 674.065 0.000 676.660 0.000
 676.660 496.905 664.245 496.905 664.245 496.035 662.715 496.035 662.715 496.905
 662.175 496.905 662.175 496.035 660.645 496.035 660.645 496.905 641.005 496.905
 641.005 496.035 639.475 496.035 639.475 496.905 638.935 496.905 638.935 496.035
 637.405 496.035 637.405 496.905 617.765 496.905 617.765 496.035 616.235 496.035
 616.235 496.905 615.695 496.905 615.695 496.035 614.165 496.035 614.165 496.905
 594.525 496.905 594.525 496.035 592.995 496.035 592.995 496.905 592.455 496.905
 592.455 496.035 590.925 496.035 590.925 496.905 571.285 496.905 571.285 496.035
 569.755 496.035 569.755 496.905 569.215 496.905 569.215 496.035 567.685 496.035
 567.685 496.905 548.045 496.905 548.045 496.035 546.515 496.035 546.515 496.905
 545.975 496.905 545.975 496.035 544.445 496.035 544.445 496.905 524.805 496.905
 524.805 496.035 523.275 496.035 523.275 496.905 522.735 496.905 522.735 496.035
 521.205 496.035 521.205 496.905 501.565 496.905 501.565 496.035 500.035 496.035
 500.035 496.905 499.495 496.905 499.495 496.035 497.965 496.035 497.965 496.905
 478.325 496.905 478.325 496.035 476.795 496.035 476.795 496.905 476.255 496.905
 476.255 496.035 474.725 496.035 474.725 496.905 455.085 496.905 455.085 496.035
 453.555 496.035 453.555 496.905 453.015 496.905 453.015 496.035 451.485 496.035
 451.485 496.905 431.845 496.905 431.845 496.035 430.315 496.035 430.315 496.905
 429.775 496.905 429.775 496.035 428.245 496.035 428.245 496.905 408.605 496.905
 408.605 496.035 407.075 496.035 407.075 496.905 406.535 496.905 406.535 496.035
 405.005 496.035 405.005 496.905 381.420 496.905 381.420 495.605 380.460 495.605
 380.460 496.905 372.015 496.905 372.015 495.605 371.055 495.605 371.055 496.905
 353.440 496.905 353.440 496.035 351.415 496.035 351.415 496.905 347.680 496.905
 347.680 496.035 345.655 496.035 345.655 496.905 341.920 496.905 341.920 496.035
 339.895 496.035 339.895 496.905 336.160 496.905 336.160 496.035 334.135 496.035
 334.135 496.905 330.400 496.905 330.400 496.035 328.375 496.035 328.375 496.905
 324.875 496.905 324.875 496.035 322.765 496.035 322.765 496.905 316.935 496.905
 316.935 496.035 314.825 496.035 314.825 496.905 308.995 496.905 308.995 496.035
 306.885 496.035 306.885 496.905 298.780 496.905 298.780 496.035 297.070 496.035
 297.070 496.905 271.655 496.905 271.655 496.035 270.125 496.035 270.125 496.905
 269.585 496.905 269.585 496.035 268.055 496.035 268.055 496.905 248.415 496.905
 248.415 496.035 246.885 496.035 246.885 496.905 246.345 496.905 246.345 496.035
 244.815 496.035 244.815 496.905 225.175 496.905 225.175 496.035 223.645 496.035
 223.645 496.905 223.105 496.905 223.105 496.035 221.575 496.035 221.575 496.905
 201.935 496.905 201.935 496.035 200.405 496.035 200.405 496.905 199.865 496.905
 199.865 496.035 198.335 496.035 198.335 496.905 178.695 496.905 178.695 496.035
 177.165 496.035 177.165 496.905 176.625 496.905 176.625 496.035 175.095 496.035
 175.095 496.905 155.455 496.905 155.455 496.035 153.925 496.035 153.925 496.905
 153.385 496.905 153.385 496.035 151.855 496.035 151.855 496.905 132.215 496.905
 132.215 496.035 130.685 496.035 130.685 496.905 130.145 496.905 130.145 496.035
 128.615 496.035 128.615 496.905 108.975 496.905 108.975 496.035 107.445 496.035
 107.445 496.905 106.905 496.905 106.905 496.035 105.375 496.035 105.375 496.905
 85.735 496.905 85.735 496.035 84.205 496.035 84.205 496.905 83.665 496.905
 83.665 496.035 82.135 496.035 82.135 496.905 62.495 496.905 62.495 496.035
 60.965 496.035 60.965 496.905 60.425 496.905 60.425 496.035 58.895 496.035
 58.895 496.905 39.255 496.905 39.255 496.035 37.725 496.035 37.725 496.905
 37.185 496.905 37.185 496.035 35.655 496.035 35.655 496.905 16.015 496.905
 16.015 496.035 14.485 496.035 14.485 496.905 13.945 496.905 13.945 496.035
 12.415 496.035 12.415 496.905 0.000 496.905 ;
LAYER METAL2 ;
POLYGON 0.000 0.000 2.545 0.000 2.545 0.920 4.175 0.920 4.175 0.000
 24.255 0.000 24.255 0.920 27.415 0.920 27.415 0.000 47.495 0.000
 47.495 0.920 50.655 0.920 50.655 0.000 70.735 0.000 70.735 0.920
 73.895 0.920 73.895 0.000 93.975 0.000 93.975 0.920 97.135 0.920
 97.135 0.000 117.215 0.000 117.215 0.920 120.375 0.920 120.375 0.000
 140.455 0.000 140.455 0.920 143.615 0.920 143.615 0.000 163.695 0.000
 163.695 0.920 166.855 0.920 166.855 0.000 186.935 0.000 186.935 0.920
 190.095 0.920 190.095 0.000 210.175 0.000 210.175 0.920 213.335 0.920
 213.335 0.000 233.415 0.000 233.415 0.920 236.575 0.920 236.575 0.000
 256.655 0.000 256.655 0.920 259.815 0.920 259.815 0.000 279.895 0.000
 279.895 0.920 281.525 0.920 281.525 0.000 296.825 0.000 296.825 1.350
 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350 307.500 1.350
 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920 325.295 0.000
 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000 335.005 0.000
 335.005 0.920 336.815 0.920 336.815 0.000 340.765 0.000 340.765 0.920
 342.575 0.920 342.575 0.000 346.525 0.000 346.525 0.920 348.335 0.920
 348.335 0.000 352.135 0.000 352.135 0.920 353.945 0.920 353.945 0.000
 360.075 0.000 360.075 0.920 361.885 0.920 361.885 0.000 368.015 0.000
 368.015 0.920 369.825 0.920 369.825 0.000 377.830 0.000 377.830 0.920
 379.640 0.920 379.640 0.000 395.135 0.000 395.135 0.920 396.765 0.920
 396.765 0.000 416.845 0.000 416.845 0.920 420.005 0.920 420.005 0.000
 440.085 0.000 440.085 0.920 443.245 0.920 443.245 0.000 463.325 0.000
 463.325 0.920 466.485 0.920 466.485 0.000 486.565 0.000 486.565 0.920
 489.725 0.920 489.725 0.000 509.805 0.000 509.805 0.920 512.965 0.920
 512.965 0.000 533.045 0.000 533.045 0.920 536.205 0.920 536.205 0.000
 556.285 0.000 556.285 0.920 559.445 0.920 559.445 0.000 579.525 0.000
 579.525 0.920 582.685 0.920 582.685 0.000 602.765 0.000 602.765 0.920
 605.925 0.920 605.925 0.000 626.005 0.000 626.005 0.920 629.165 0.920
 629.165 0.000 649.245 0.000 649.245 0.920 652.405 0.920 652.405 0.000
 672.485 0.000 672.485 0.920 674.115 0.920 674.115 0.000 676.660 0.000
 676.660 496.905 664.295 496.905 664.295 495.985 662.665 495.985 662.665 496.905
 662.225 496.905 662.225 495.985 660.595 495.985 660.595 496.905 641.055 496.905
 641.055 495.985 639.425 495.985 639.425 496.905 638.985 496.905 638.985 495.985
 637.355 495.985 637.355 496.905 617.815 496.905 617.815 495.985 616.185 495.985
 616.185 496.905 615.745 496.905 615.745 495.985 614.115 495.985 614.115 496.905
 594.575 496.905 594.575 495.985 592.945 495.985 592.945 496.905 592.505 496.905
 592.505 495.985 590.875 495.985 590.875 496.905 571.335 496.905 571.335 495.985
 569.705 495.985 569.705 496.905 569.265 496.905 569.265 495.985 567.635 495.985
 567.635 496.905 548.095 496.905 548.095 495.985 546.465 495.985 546.465 496.905
 546.025 496.905 546.025 495.985 544.395 495.985 544.395 496.905 524.855 496.905
 524.855 495.985 523.225 495.985 523.225 496.905 522.785 496.905 522.785 495.985
 521.155 495.985 521.155 496.905 501.615 496.905 501.615 495.985 499.985 495.985
 499.985 496.905 499.545 496.905 499.545 495.985 497.915 495.985 497.915 496.905
 478.375 496.905 478.375 495.985 476.745 495.985 476.745 496.905 476.305 496.905
 476.305 495.985 474.675 495.985 474.675 496.905 455.135 496.905 455.135 495.985
 453.505 495.985 453.505 496.905 453.065 496.905 453.065 495.985 451.435 495.985
 451.435 496.905 431.895 496.905 431.895 495.985 430.265 495.985 430.265 496.905
 429.825 496.905 429.825 495.985 428.195 495.985 428.195 496.905 408.655 496.905
 408.655 495.985 407.025 495.985 407.025 496.905 406.585 496.905 406.585 495.985
 404.955 495.985 404.955 496.905 381.470 496.905 381.470 495.555 380.410 495.555
 380.410 496.905 372.065 496.905 372.065 495.555 371.005 495.555 371.005 496.905
 353.175 496.905 353.175 495.985 351.365 495.985 351.365 496.905 347.415 496.905
 347.415 495.985 345.605 495.985 345.605 496.905 341.655 496.905 341.655 495.985
 339.845 495.985 339.845 496.905 335.895 496.905 335.895 495.985 334.085 495.985
 334.085 496.905 330.135 496.905 330.135 495.985 328.325 495.985 328.325 496.905
 324.525 496.905 324.525 495.985 322.715 495.985 322.715 496.905 316.585 496.905
 316.585 495.985 314.775 495.985 314.775 496.905 308.645 496.905 308.645 495.985
 306.835 495.985 306.835 496.905 298.830 496.905 298.830 495.985 297.020 495.985
 297.020 496.905 271.705 496.905 271.705 495.985 270.075 495.985 270.075 496.905
 269.635 496.905 269.635 495.985 268.005 495.985 268.005 496.905 248.465 496.905
 248.465 495.985 246.835 495.985 246.835 496.905 246.395 496.905 246.395 495.985
 244.765 495.985 244.765 496.905 225.225 496.905 225.225 495.985 223.595 495.985
 223.595 496.905 223.155 496.905 223.155 495.985 221.525 495.985 221.525 496.905
 201.985 496.905 201.985 495.985 200.355 495.985 200.355 496.905 199.915 496.905
 199.915 495.985 198.285 495.985 198.285 496.905 178.745 496.905 178.745 495.985
 177.115 495.985 177.115 496.905 176.675 496.905 176.675 495.985 175.045 495.985
 175.045 496.905 155.505 496.905 155.505 495.985 153.875 495.985 153.875 496.905
 153.435 496.905 153.435 495.985 151.805 495.985 151.805 496.905 132.265 496.905
 132.265 495.985 130.635 495.985 130.635 496.905 130.195 496.905 130.195 495.985
 128.565 495.985 128.565 496.905 109.025 496.905 109.025 495.985 107.395 495.985
 107.395 496.905 106.955 496.905 106.955 495.985 105.325 495.985 105.325 496.905
 85.785 496.905 85.785 495.985 84.155 495.985 84.155 496.905 83.715 496.905
 83.715 495.985 82.085 495.985 82.085 496.905 62.545 496.905 62.545 495.985
 60.915 495.985 60.915 496.905 60.475 496.905 60.475 495.985 58.845 495.985
 58.845 496.905 39.305 496.905 39.305 495.985 37.675 495.985 37.675 496.905
 37.235 496.905 37.235 495.985 35.605 495.985 35.605 496.905 16.065 496.905
 16.065 495.985 14.435 495.985 14.435 496.905 13.995 496.905 13.995 495.985
 12.365 495.985 12.365 496.905 0.000 496.905 ;
LAYER METAL3 ;
POLYGON 0.000 0.000 2.545 0.000 2.545 0.920 4.175 0.920 4.175 0.000
 24.255 0.000 24.255 0.920 27.415 0.920 27.415 0.000 47.495 0.000
 47.495 0.920 50.655 0.920 50.655 0.000 70.735 0.000 70.735 0.920
 73.895 0.920 73.895 0.000 93.975 0.000 93.975 0.920 97.135 0.920
 97.135 0.000 117.215 0.000 117.215 0.920 120.375 0.920 120.375 0.000
 140.455 0.000 140.455 0.920 143.615 0.920 143.615 0.000 163.695 0.000
 163.695 0.920 166.855 0.920 166.855 0.000 186.935 0.000 186.935 0.920
 190.095 0.920 190.095 0.000 210.175 0.000 210.175 0.920 213.335 0.920
 213.335 0.000 233.415 0.000 233.415 0.920 236.575 0.920 236.575 0.000
 256.655 0.000 256.655 0.920 259.815 0.920 259.815 0.000 279.895 0.000
 279.895 0.920 281.525 0.920 281.525 0.000 296.825 0.000 296.825 1.350
 297.885 1.350 297.885 0.000 306.440 0.000 306.440 1.350 307.500 1.350
 307.500 0.000 323.485 0.000 323.485 0.920 325.295 0.920 325.295 0.000
 329.245 0.000 329.245 0.920 331.055 0.920 331.055 0.000 335.005 0.000
 335.005 0.920 336.815 0.920 336.815 0.000 340.765 0.000 340.765 0.920
 342.575 0.920 342.575 0.000 346.525 0.000 346.525 0.920 348.335 0.920
 348.335 0.000 352.135 0.000 352.135 0.920 353.945 0.920 353.945 0.000
 360.075 0.000 360.075 0.920 361.885 0.920 361.885 0.000 368.015 0.000
 368.015 0.920 369.825 0.920 369.825 0.000 377.830 0.000 377.830 0.920
 379.640 0.920 379.640 0.000 395.135 0.000 395.135 0.920 396.765 0.920
 396.765 0.000 416.845 0.000 416.845 0.920 420.005 0.920 420.005 0.000
 440.085 0.000 440.085 0.920 443.245 0.920 443.245 0.000 463.325 0.000
 463.325 0.920 466.485 0.920 466.485 0.000 486.565 0.000 486.565 0.920
 489.725 0.920 489.725 0.000 509.805 0.000 509.805 0.920 512.965 0.920
 512.965 0.000 533.045 0.000 533.045 0.920 536.205 0.920 536.205 0.000
 556.285 0.000 556.285 0.920 559.445 0.920 559.445 0.000 579.525 0.000
 579.525 0.920 582.685 0.920 582.685 0.000 602.765 0.000 602.765 0.920
 605.925 0.920 605.925 0.000 626.005 0.000 626.005 0.920 629.165 0.920
 629.165 0.000 649.245 0.000 649.245 0.920 652.405 0.920 652.405 0.000
 672.485 0.000 672.485 0.920 674.115 0.920 674.115 0.000 676.660 0.000
 676.660 496.905 664.295 496.905 664.295 495.985 662.665 495.985 662.665 496.905
 662.225 496.905 662.225 495.985 660.595 495.985 660.595 496.905 641.055 496.905
 641.055 495.985 639.425 495.985 639.425 496.905 638.985 496.905 638.985 495.985
 637.355 495.985 637.355 496.905 617.815 496.905 617.815 495.985 616.185 495.985
 616.185 496.905 615.745 496.905 615.745 495.985 614.115 495.985 614.115 496.905
 594.575 496.905 594.575 495.985 592.945 495.985 592.945 496.905 592.505 496.905
 592.505 495.985 590.875 495.985 590.875 496.905 571.335 496.905 571.335 495.985
 569.705 495.985 569.705 496.905 569.265 496.905 569.265 495.985 567.635 495.985
 567.635 496.905 548.095 496.905 548.095 495.985 546.465 495.985 546.465 496.905
 546.025 496.905 546.025 495.985 544.395 495.985 544.395 496.905 524.855 496.905
 524.855 495.985 523.225 495.985 523.225 496.905 522.785 496.905 522.785 495.985
 521.155 495.985 521.155 496.905 501.615 496.905 501.615 495.985 499.985 495.985
 499.985 496.905 499.545 496.905 499.545 495.985 497.915 495.985 497.915 496.905
 478.375 496.905 478.375 495.985 476.745 495.985 476.745 496.905 476.305 496.905
 476.305 495.985 474.675 495.985 474.675 496.905 455.135 496.905 455.135 495.985
 453.505 495.985 453.505 496.905 453.065 496.905 453.065 495.985 451.435 495.985
 451.435 496.905 431.895 496.905 431.895 495.985 430.265 495.985 430.265 496.905
 429.825 496.905 429.825 495.985 428.195 495.985 428.195 496.905 408.655 496.905
 408.655 495.985 407.025 495.985 407.025 496.905 406.585 496.905 406.585 495.985
 404.955 495.985 404.955 496.905 381.470 496.905 381.470 495.555 380.410 495.555
 380.410 496.905 372.065 496.905 372.065 495.555 371.005 495.555 371.005 496.905
 353.175 496.905 353.175 495.985 351.365 495.985 351.365 496.905 347.415 496.905
 347.415 495.985 345.605 495.985 345.605 496.905 341.655 496.905 341.655 495.985
 339.845 495.985 339.845 496.905 335.895 496.905 335.895 495.985 334.085 495.985
 334.085 496.905 330.135 496.905 330.135 495.985 328.325 495.985 328.325 496.905
 324.525 496.905 324.525 495.985 322.715 495.985 322.715 496.905 316.585 496.905
 316.585 495.985 314.775 495.985 314.775 496.905 308.645 496.905 308.645 495.985
 306.835 495.985 306.835 496.905 298.830 496.905 298.830 495.985 297.020 495.985
 297.020 496.905 271.705 496.905 271.705 495.985 270.075 495.985 270.075 496.905
 269.635 496.905 269.635 495.985 268.005 495.985 268.005 496.905 248.465 496.905
 248.465 495.985 246.835 495.985 246.835 496.905 246.395 496.905 246.395 495.985
 244.765 495.985 244.765 496.905 225.225 496.905 225.225 495.985 223.595 495.985
 223.595 496.905 223.155 496.905 223.155 495.985 221.525 495.985 221.525 496.905
 201.985 496.905 201.985 495.985 200.355 495.985 200.355 496.905 199.915 496.905
 199.915 495.985 198.285 495.985 198.285 496.905 178.745 496.905 178.745 495.985
 177.115 495.985 177.115 496.905 176.675 496.905 176.675 495.985 175.045 495.985
 175.045 496.905 155.505 496.905 155.505 495.985 153.875 495.985 153.875 496.905
 153.435 496.905 153.435 495.985 151.805 495.985 151.805 496.905 132.265 496.905
 132.265 495.985 130.635 495.985 130.635 496.905 130.195 496.905 130.195 495.985
 128.565 495.985 128.565 496.905 109.025 496.905 109.025 495.985 107.395 495.985
 107.395 496.905 106.955 496.905 106.955 495.985 105.325 495.985 105.325 496.905
 85.785 496.905 85.785 495.985 84.155 495.985 84.155 496.905 83.715 496.905
 83.715 495.985 82.085 495.985 82.085 496.905 62.545 496.905 62.545 495.985
 60.915 495.985 60.915 496.905 60.475 496.905 60.475 495.985 58.845 495.985
 58.845 496.905 39.305 496.905 39.305 495.985 37.675 495.985 37.675 496.905
 37.235 496.905 37.235 495.985 35.605 495.985 35.605 496.905 16.065 496.905
 16.065 495.985 14.435 495.985 14.435 496.905 13.995 496.905 13.995 495.985
 12.365 495.985 12.365 496.905 0.000 496.905 ;
END
END FRAM512
END LIBRARY
